netcdf tmp_xarrayanon {
dimensions:
	_Anonymous_Dim_2 = 2 ;
	_Anonymous_Dim_3 = 3 ;
variables:
 	int i(_Anonymous_Dim_2, _Anonymous_Dim_3) ;
data:

 i =
  _, _, _,
  _, _, _ ;
}
