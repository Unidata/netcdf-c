[0] /.nczarr : (0) ||
