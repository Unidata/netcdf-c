netcdf t_ncgen {
dimensions:
	dim1 = 1 ;
variables:
	int var1 ;
}
