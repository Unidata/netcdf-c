netcdf y {
dimensions:
	Dr = UNLIMITED ; // (2 currently)
	D1 = 1 ;
	D2 = 2 ;
	D3 = 3 ;
        U=unlimited;
variables:
 char cuu(Dr,D2,U);
data:
 cuu = {{"a","def"}}, {{"xy"}};

}
