testmap.nzf
testmap.nzf/.nczarr : ||
