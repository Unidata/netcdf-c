netcdf tim {
types:
  byte enum e1{pass=0, fail=1, undefined=2};
  byte enum e2{defined=0, undefined=1};
variables:
  e1 test1;
  e2 test2;
  e2 test3;
data:
  test1=pass;
  test2=e1.undefined;
  test3=/e1.fail;
} 
