netcdf tmp_purezarr {
dimensions:
	x = 2 ;
	y = 5 ;
variables:
	int i(x, y) ;
data:

 i =
  _, _, _, _, _,
  _, _, _, _, _ ;
}
