netcdf ref_oldformat {
dimensions:
	lat = 8 ;
	_zdim_8 = 8 ;
	_zdim_10 = 10 ;
variables:
	int lat(lat) ;
		lat:_FillValue = -1 ;
		string lat:lat_attr = "latitude" ;
data:

 lat = 1, 2, 3, 4, 5, 6, 7, 8 ;

group: g1 {
  variables:
  	int pos(_zdim_8, _zdim_10) ;
  		pos:_FillValue = -1 ;
  		string pos:pos_attr = "latXlon" ;

  // group attributes:
  		:g1_attr = 17 ;
  data:

   pos =
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _ ;
  } // group g1
}
