netcdf c0 {
dimensions:
	Dr = UNLIMITED ;
	D1 = 1 ;
	D2 = 2 ;
	D3 = 3 ;
variables:
  char c;
  car c1(D1);
  char c13(D1, D3) ;
  char c31(D3, D1) ;
  char c111(D1, D1, D1) ;
  char c123(D1, D2, D3) ;
  char c213(D2, D1, D3) ;
  char c231(D2, D3, D1) ;
  char cr(Dr) ;
  char cra(Dr) ;
  char c2a(D2) ;
  char cr1(Dr, D1) ;
  char cr2(Dr, D2) ;
  char cr21(Dr, D2, D1) ;
  char cr33(Dr, D3, D3) ;
data:
  c = "2" ;
  c1 = "";
  c2 = "a", "b" ;
  c2a = 'a', 'b' ;
  c3 = "\001\300." ;
  c13 = "\tb\177" ;
  c31 = "+", "-", " " ;
  c111 = "@" ;
  c123 = "one", "2" ;
  c213 = "1", "two" ;
  c231 = "@", "D", "H", "H", "L", "P" ;
  cra = "ab" ;
  cr = "a","b" ;
  cr2 =  "@",  "D",  "H",  "L" ;
  cr21 =  "@",  "D",  "H",  "L" ;
  cr33 =  "1", "two",  "3",  "4",  "5",  "six" ;
}
 
