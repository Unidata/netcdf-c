netcdf ref_tst_perdimspecs {
dimensions:
	lon = 40 ;
	lat = 41 ;
	time = 42;
variables:
	float lon(lon) ;
	float lat(lat) ;
	double time(time) ;
	float tas(time, lat, lon) ;
}
