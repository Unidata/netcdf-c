netcdf ref_oldformat {
dimensions:
	lat = 8 ;
variables:
	int lat(lat) ;
		lat:_FillValue = -1 ;
		lat:lat_attr = "latitude" ;
data:

 lat = 1, 2, 3, 4, 5, 6, 7, 8 ;

group: g1 {
  dimensions:
  	lon = 10 ;
  variables:
  	int pos(lat, lon) ;
  		pos:_FillValue = -1 ;
  		pos:pos_attr = "latXlon" ;

  // group attributes:
  		:g1_attr = 17 ;
  data:

   pos =
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _ ;
  } // group g1
}
