netcdf test_corrupt_magic {
dimensions:
	recNum = 8;
variables:
	string UTC_time(recNum) ;
data:

 UTC_time = "2012-03-04 03:54:19", "2012-03-04 03:54:42", 
    "2012-03-04 03:54:59", "2012-03-04 03:55:20", "2012-03-04 03:55:43", 
    "2012-03-04 03:56:09", "2012-03-04 03:56:41", "2012-03-04 03:57:12" ;
}
