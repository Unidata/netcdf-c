netcdf type_ancestor_subgroup {
types:
  ubyte enum test_enum_type {OPTION1 = 0, OPTION2 = 1, OPTION3 = 2} ;

group: test_group {
  variables:
  	test_enum_type test_variable ;
  		test_enum_type test_variable:_FillValue = OPTION1 ;
  group: sub_group {
      types:
      ubyte enum test_enum_type {OPTION1 = 0, OPTION2 = 1, OPTION3 = 2} ;
  } // group sub_group

  } // group test_group
}
