netcdf testmap {

group: _nczarr {
  } // group _nczarr
}
