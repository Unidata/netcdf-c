netcdf OR_ABI-L1b-RadF-M6C01_G16_s20220011800205_e20220011809513_c20220011809562 {
dimensions:
	y = 10848 ;
	x = 10848 ;
	number_of_time_bounds = 2 ;
	band = 1 ;
	number_of_image_bounds = 2 ;
	num_star_looks = 24 ;
variables:
	short Rad(y, x) ;
		Rad:_FillValue = 1023s ;
		Rad:long_name = "ABI L1b Radiances" ;
		Rad:standard_name = "toa_outgoing_radiance_per_unit_wavelength" ;
		Rad:_Unsigned = "true" ;
		Rad:sensor_band_bit_depth = 10b ;
		Rad:valid_range = 0s, 1022s ;
		Rad:scale_factor = 0.8121064f ;
		Rad:add_offset = -25.93665f ;
		Rad:units = "W m-2 sr-1 um-1" ;
		Rad:resolution = "y: 0.000028 rad x: 0.000028 rad" ;
		Rad:coordinates = "band_id band_wavelength t y x" ;
		Rad:grid_mapping = "goes_imager_projection" ;
		Rad:cell_methods = "t: point area: point" ;
		Rad:ancillary_variables = "DQF" ;
	byte DQF(y, x) ;
		DQF:_FillValue = -1b ;
		DQF:long_name = "ABI L1b Radiances data quality flags" ;
		DQF:standard_name = "status_flag" ;
		DQF:_Unsigned = "true" ;
		DQF:valid_range = 0b, 4b ;
		DQF:units = "1" ;
		DQF:coordinates = "band_id band_wavelength t y x" ;
		DQF:grid_mapping = "goes_imager_projection" ;
		DQF:cell_methods = "t: point area: point" ;
		DQF:flag_values = 0b, 1b, 2b, 3b, 4b ;
		DQF:flag_meanings = "good_pixel_qf conditionally_usable_pixel_qf out_of_range_pixel_qf no_value_pixel_qf focal_plane_temperature_threshold_exceeded_qf" ;
		DQF:number_of_qf_values = 5b ;
		DQF:percent_good_pixel_qf = 0.998999f ;
		DQF:percent_conditionally_usable_pixel_qf = 5.e-07f ;
		DQF:percent_out_of_range_pixel_qf = 0.0009925f ;
		DQF:percent_no_value_pixel_qf = 8.e-06f ;
		DQF:percent_focal_plane_temperature_threshold_exceeded_qf = 0.f ;
	double t ;
		t:long_name = "J2000 epoch mid-point between the start and end image scan in seconds" ;
		t:standard_name = "time" ;
		t:units = "seconds since 2000-01-01 12:00:00" ;
		t:axis = "T" ;
		t:bounds = "time_bounds" ;
	short y(y) ;
		y:scale_factor = -2.8e-05f ;
		y:add_offset = 0.151858f ;
		y:units = "rad" ;
		y:axis = "Y" ;
		y:long_name = "GOES fixed grid projection y-coordinate" ;
		y:standard_name = "projection_y_coordinate" ;
	short x(x) ;
		x:scale_factor = 2.8e-05f ;
		x:add_offset = -0.151858f ;
		x:units = "rad" ;
		x:axis = "X" ;
		x:long_name = "GOES fixed grid projection x-coordinate" ;
		x:standard_name = "projection_x_coordinate" ;
	double time_bounds(number_of_time_bounds) ;
		time_bounds:long_name = "Scan start and end times in seconds since epoch (2000-01-01 12:00:00)" ;
	int goes_imager_projection ;
		goes_imager_projection:long_name = "GOES-R ABI fixed grid projection" ;
		goes_imager_projection:grid_mapping_name = "geostationary" ;
		goes_imager_projection:perspective_point_height = 35786023. ;
		goes_imager_projection:semi_major_axis = 6378137. ;
		goes_imager_projection:semi_minor_axis = 6356752.31414 ;
		goes_imager_projection:inverse_flattening = 298.2572221 ;
		goes_imager_projection:latitude_of_projection_origin = 0. ;
		goes_imager_projection:longitude_of_projection_origin = -75. ;
		goes_imager_projection:sweep_angle_axis = "x" ;
	float y_image ;
		y_image:long_name = "GOES-R fixed grid projection y-coordinate center of image" ;
		y_image:standard_name = "projection_y_coordinate" ;
		y_image:units = "rad" ;
		y_image:axis = "Y" ;
	float y_image_bounds(number_of_image_bounds) ;
		y_image_bounds:long_name = "GOES-R fixed grid projection y-coordinate north/south extent of image" ;
		y_image_bounds:units = "rad" ;
	float x_image ;
		x_image:long_name = "GOES-R fixed grid projection x-coordinate center of image" ;
		x_image:standard_name = "projection_x_coordinate" ;
		x_image:units = "rad" ;
		x_image:axis = "X" ;
	float x_image_bounds(number_of_image_bounds) ;
		x_image_bounds:long_name = "GOES-R fixed grid projection x-coordinate west/east extent of image" ;
		x_image_bounds:units = "rad" ;
	float nominal_satellite_subpoint_lat ;
		nominal_satellite_subpoint_lat:long_name = "nominal satellite subpoint latitude (platform latitude)" ;
		nominal_satellite_subpoint_lat:standard_name = "latitude" ;
		nominal_satellite_subpoint_lat:_FillValue = -999.f ;
		nominal_satellite_subpoint_lat:units = "degrees_north" ;
	float nominal_satellite_subpoint_lon ;
		nominal_satellite_subpoint_lon:long_name = "nominal satellite subpoint longitude (platform longitude)" ;
		nominal_satellite_subpoint_lon:standard_name = "longitude" ;
		nominal_satellite_subpoint_lon:_FillValue = -999.f ;
		nominal_satellite_subpoint_lon:units = "degrees_east" ;
	float nominal_satellite_height ;
		nominal_satellite_height:long_name = "nominal satellite height above GRS 80 ellipsoid (platform altitude)" ;
		nominal_satellite_height:standard_name = "height_above_reference_ellipsoid" ;
		nominal_satellite_height:_FillValue = -999.f ;
		nominal_satellite_height:units = "km" ;
	float geospatial_lat_lon_extent ;
		geospatial_lat_lon_extent:long_name = "geospatial latitude and longitude references" ;
		geospatial_lat_lon_extent:geospatial_westbound_longitude = -156.2995f ;
		geospatial_lat_lon_extent:geospatial_northbound_latitude = 81.3282f ;
		geospatial_lat_lon_extent:geospatial_eastbound_longitude = 6.2995f ;
		geospatial_lat_lon_extent:geospatial_southbound_latitude = -81.3282f ;
		geospatial_lat_lon_extent:geospatial_lat_center = 0.f ;
		geospatial_lat_lon_extent:geospatial_lon_center = -75.f ;
		geospatial_lat_lon_extent:geospatial_lat_nadir = 0.f ;
		geospatial_lat_lon_extent:geospatial_lon_nadir = -75.f ;
		geospatial_lat_lon_extent:geospatial_lat_units = "degrees_north" ;
		geospatial_lat_lon_extent:geospatial_lon_units = "degrees_east" ;
	byte yaw_flip_flag ;
		yaw_flip_flag:long_name = "Flag indicating the spacecraft is operating in yaw flip configuration" ;
		yaw_flip_flag:_Unsigned = "true" ;
		yaw_flip_flag:_FillValue = -1b ;
		yaw_flip_flag:valid_range = 0b, 1b ;
		yaw_flip_flag:units = "1" ;
		yaw_flip_flag:coordinates = "t" ;
		yaw_flip_flag:flag_values = 0b, 1b ;
		yaw_flip_flag:flag_meanings = "false true" ;
	byte band_id(band) ;
		band_id:long_name = "ABI band number" ;
		band_id:standard_name = "sensor_band_identifier" ;
		band_id:units = "1" ;
	float band_wavelength(band) ;
		band_wavelength:long_name = "ABI band central wavelength" ;
		band_wavelength:standard_name = "sensor_band_central_radiation_wavelength" ;
		band_wavelength:units = "um" ;
	float esun ;
		esun:long_name = "bandpass-weighted solar irradiance at the mean Earth-Sun distance" ;
		esun:standard_name = "toa_shortwave_irradiance_per_unit_wavelength" ;
		esun:_FillValue = -999.f ;
		esun:units = "W m-2 um-1" ;
		esun:coordinates = "band_id band_wavelength t" ;
		esun:cell_methods = "t: mean" ;
	float kappa0 ;
		kappa0:long_name = "Inverse of the incoming top of atmosphere radiance at current earth-sun distance (PI d2 esun-1)-1, where d is the ratio of instantaneous Earth-Sun distance divided by the mean Earth-Sun distance, esun is the bandpass-weighted solar irradiance and PI is a standard constant used to convert ABI L1b radiance to reflectance" ;
		kappa0:_FillValue = -999.f ;
		kappa0:units = "(W m-2 um-1)-1" ;
		kappa0:coordinates = "band_id band_wavelength t" ;
		kappa0:cell_methods = "t: mean" ;
	float planck_fk1 ;
		planck_fk1:long_name = "wavenumber-dependent coefficient (2 h c2/ nu3) used in the ABI emissive band monochromatic brightness temperature computation, where nu =central wavenumber and h and c are standard constants" ;
		planck_fk1:_FillValue = -999.f ;
		planck_fk1:units = "W m-1" ;
		planck_fk1:coordinates = "band_id band_wavelength" ;
	float planck_fk2 ;
		planck_fk2:long_name = "wavenumber-dependent coefficient (h c nu/b) used in the ABI emissive band monochromatic brightness temperature computation, where nu = central wavenumber and h, c, and b are standard constants" ;
		planck_fk2:_FillValue = -999.f ;
		planck_fk2:units = "K" ;
		planck_fk2:coordinates = "band_id band_wavelength" ;
	float planck_bc1 ;
		planck_bc1:long_name = "spectral bandpass correction offset for brightness temperature (B(nu) - bc_1)/bc_2 where B()=planck_function() and nu=wavenumber" ;
		planck_bc1:_FillValue = -999.f ;
		planck_bc1:units = "K" ;
		planck_bc1:coordinates = "band_id band_wavelength" ;
	float planck_bc2 ;
		planck_bc2:long_name = "spectral bandpass correction scale factor for brightness temperature (B(nu) - bc_1)/bc_2 where B()=planck_function() and nu=wavenumber" ;
		planck_bc2:_FillValue = -999.f ;
		planck_bc2:units = "1" ;
		planck_bc2:coordinates = "band_id band_wavelength" ;
	int valid_pixel_count ;
		valid_pixel_count:long_name = "number of good and conditionally usable pixels" ;
		valid_pixel_count:_FillValue = -1 ;
		valid_pixel_count:units = "count" ;
		valid_pixel_count:coordinates = "band_id band_wavelength t y_image x_image" ;
		valid_pixel_count:grid_mapping = "goes_imager_projection" ;
		valid_pixel_count:cell_methods = "t: sum area: sum (interval: 0.000028 rad comment: good and conditionally usable quality pixels only)" ;
	int missing_pixel_count ;
		missing_pixel_count:long_name = "number of missing pixels" ;
		missing_pixel_count:_FillValue = -1 ;
		missing_pixel_count:units = "count" ;
		missing_pixel_count:coordinates = "band_id band_wavelength t y_image x_image" ;
		missing_pixel_count:grid_mapping = "goes_imager_projection" ;
		missing_pixel_count:cell_methods = "t: sum area: sum (interval: 0.000028 rad comment: missing ABI fixed grid pixels only)" ;
	int saturated_pixel_count ;
		saturated_pixel_count:long_name = "number of saturated pixels" ;
		saturated_pixel_count:_FillValue = -1 ;
		saturated_pixel_count:units = "count" ;
		saturated_pixel_count:coordinates = "band_id band_wavelength t y_image x_image" ;
		saturated_pixel_count:grid_mapping = "goes_imager_projection" ;
		saturated_pixel_count:cell_methods = "t: sum area: sum (interval: 0.000028 rad comment: radiometrically saturated geolocated/not missing pixels only)" ;
	int undersaturated_pixel_count ;
		undersaturated_pixel_count:long_name = "number of undersaturated pixels" ;
		undersaturated_pixel_count:_FillValue = -1 ;
		undersaturated_pixel_count:units = "count" ;
		undersaturated_pixel_count:coordinates = "band_id band_wavelength t y_image x_image" ;
		undersaturated_pixel_count:grid_mapping = "goes_imager_projection" ;
		undersaturated_pixel_count:cell_methods = "t: sum area: sum (interval: 0.000028 rad comment: radiometrically undersaturated geolocated/not missing pixels only)" ;
	int focal_plane_temperature_threshold_exceeded_count ;
		focal_plane_temperature_threshold_exceeded_count:long_name = "number of pixels whose temperatures exceeded the threshold" ;
		focal_plane_temperature_threshold_exceeded_count:_FillValue = -1 ;
		focal_plane_temperature_threshold_exceeded_count:units = "count" ;
		focal_plane_temperature_threshold_exceeded_count:coordinates = "band_id band_wavelength t y_image x_image" ;
		focal_plane_temperature_threshold_exceeded_count:grid_mapping = "goes_imager_projection" ;
		focal_plane_temperature_threshold_exceeded_count:cell_methods = "t: sum area: sum (interval: 0.000028 rad comment: temperature exceeded pixels only)" ;
	float min_radiance_value_of_valid_pixels ;
		min_radiance_value_of_valid_pixels:long_name = "minimum radiance value of pixels" ;
		min_radiance_value_of_valid_pixels:standard_name = "toa_outgoing_radiance_per_unit_wavelength" ;
		min_radiance_value_of_valid_pixels:_FillValue = -999.f ;
		min_radiance_value_of_valid_pixels:valid_range = -25.93665f, 804.0361f ;
		min_radiance_value_of_valid_pixels:units = "W m-2 sr-1 um-1" ;
		min_radiance_value_of_valid_pixels:coordinates = "band_id band_wavelength t y_image x_image" ;
		min_radiance_value_of_valid_pixels:grid_mapping = "goes_imager_projection" ;
		min_radiance_value_of_valid_pixels:cell_methods = "t: sum area: minimum (interval: 0.000028 rad comment: good and conditionally usable quality pixels only)" ;
	float max_radiance_value_of_valid_pixels ;
		max_radiance_value_of_valid_pixels:long_name = "maximum radiance value of pixels" ;
		max_radiance_value_of_valid_pixels:standard_name = "toa_outgoing_radiance_per_unit_wavelength" ;
		max_radiance_value_of_valid_pixels:_FillValue = -999.f ;
		max_radiance_value_of_valid_pixels:valid_range = -25.93665f, 804.0361f ;
		max_radiance_value_of_valid_pixels:units = "W m-2 sr-1 um-1" ;
		max_radiance_value_of_valid_pixels:coordinates = "band_id band_wavelength t y_image x_image" ;
		max_radiance_value_of_valid_pixels:grid_mapping = "goes_imager_projection" ;
		max_radiance_value_of_valid_pixels:cell_methods = "t: sum area: maximum (interval: 0.000028 rad comment: good and conditionally usable quality pixels only)" ;
	float mean_radiance_value_of_valid_pixels ;
		mean_radiance_value_of_valid_pixels:long_name = "mean radiance value of pixels" ;
		mean_radiance_value_of_valid_pixels:standard_name = "toa_outgoing_radiance_per_unit_wavelength" ;
		mean_radiance_value_of_valid_pixels:_FillValue = -999.f ;
		mean_radiance_value_of_valid_pixels:valid_range = -25.93665f, 804.0361f ;
		mean_radiance_value_of_valid_pixels:units = "W m-2 sr-1 um-1" ;
		mean_radiance_value_of_valid_pixels:coordinates = "band_id band_wavelength t y_image x_image" ;
		mean_radiance_value_of_valid_pixels:grid_mapping = "goes_imager_projection" ;
		mean_radiance_value_of_valid_pixels:cell_methods = "t: sum area: mean (interval: 0.000028 rad comment: good and conditionally usable quality pixels only)" ;
	float std_dev_radiance_value_of_valid_pixels ;
		std_dev_radiance_value_of_valid_pixels:long_name = "standard deviation of radiance values of pixels" ;
		std_dev_radiance_value_of_valid_pixels:standard_name = "toa_outgoing_radiance_per_unit_wavelength" ;
		std_dev_radiance_value_of_valid_pixels:_FillValue = -999.f ;
		std_dev_radiance_value_of_valid_pixels:units = "W m-2 sr-1 um-1" ;
		std_dev_radiance_value_of_valid_pixels:coordinates = "band_id band_wavelength t y_image x_image" ;
		std_dev_radiance_value_of_valid_pixels:grid_mapping = "goes_imager_projection" ;
		std_dev_radiance_value_of_valid_pixels:cell_methods = "t: sum area: standard_deviation (interval: 0.000028 rad comment: good and conditionally usable quality pixels only)" ;
	float maximum_focal_plane_temperature ;
		maximum_focal_plane_temperature:long_name = "maximum focal plane temperature value" ;
		maximum_focal_plane_temperature:_FillValue = -999.f ;
		maximum_focal_plane_temperature:valid_range = 0.f, 999.f ;
		maximum_focal_plane_temperature:units = "K" ;
	float focal_plane_temperature_threshold_increasing ;
		focal_plane_temperature_threshold_increasing:long_name = "focal plane temperature threshold increasing bounds value" ;
		focal_plane_temperature_threshold_increasing:_FillValue = -999.f ;
		focal_plane_temperature_threshold_increasing:valid_range = 0.f, 999.f ;
		focal_plane_temperature_threshold_increasing:units = "K" ;
	float focal_plane_temperature_threshold_decreasing ;
		focal_plane_temperature_threshold_decreasing:long_name = "focal plane temperature threshold decreasing bounds value" ;
		focal_plane_temperature_threshold_decreasing:_FillValue = -999.f ;
		focal_plane_temperature_threshold_decreasing:valid_range = 0.f, 999.f ;
		focal_plane_temperature_threshold_decreasing:units = "K" ;
	float percent_uncorrectable_L0_errors ;
		percent_uncorrectable_L0_errors:long_name = "percent data lost due to uncorrectable L0 errors" ;
		percent_uncorrectable_L0_errors:_FillValue = -999.f ;
		percent_uncorrectable_L0_errors:valid_range = 0.f, 1.f ;
		percent_uncorrectable_L0_errors:units = "percent" ;
		percent_uncorrectable_L0_errors:coordinates = "t y_image x_image" ;
		percent_uncorrectable_L0_errors:grid_mapping = "goes_imager_projection" ;
		percent_uncorrectable_L0_errors:cell_methods = "t: sum area: sum (uncorrectable L0 errors only)" ;
	float earth_sun_distance_anomaly_in_AU ;
		earth_sun_distance_anomaly_in_AU:long_name = "earth sun distance anomaly in astronomical units" ;
		earth_sun_distance_anomaly_in_AU:_FillValue = -999.f ;
		earth_sun_distance_anomaly_in_AU:units = "ua" ;
		earth_sun_distance_anomaly_in_AU:coordinates = "t" ;
		earth_sun_distance_anomaly_in_AU:cell_methods = "t: mean" ;
	int algorithm_dynamic_input_data_container ;
		algorithm_dynamic_input_data_container:long_name = "container for filenames of dynamic algorithm input data" ;
		algorithm_dynamic_input_data_container:input_ABI_L0_data = "OR_ABI-L0-F-M6_G16_s20220011800205_e20220011809513_c*.nc" ;
	int processing_parm_version_container ;
		processing_parm_version_container:long_name = "container for processing parameter filenames" ;
		processing_parm_version_container:L1b_processing_parm_version = "OR-PARM-RAD_G16_v01r00.zip" ;
	int algorithm_product_version_container ;
		algorithm_product_version_container:long_name = "container for algorithm package filename and product version" ;
		algorithm_product_version_container:algorithm_version = "OR_ABI-L1b-ALG-RAD_v01r00.zip" ;
		algorithm_product_version_container:product_version = "v01r00" ;
	double t_star_look(num_star_looks) ;
		t_star_look:long_name = "J2000 epoch time of star observed in seconds" ;
		t_star_look:standard_name = "time" ;
		t_star_look:units = "seconds since 2000-01-01 12:00:00" ;
		t_star_look:axis = "T" ;
	float band_wavelength_star_look(num_star_looks) ;
		band_wavelength_star_look:long_name = "ABI band central wavelength associated with observed star" ;
		band_wavelength_star_look:standard_name = "sensor_band_central_radiation_wavelength" ;
		band_wavelength_star_look:units = "um" ;
	short star_id(num_star_looks) ;
		star_id:long_name = "ABI star catalog identifier associated with observed star" ;
		star_id:_Unsigned = "true" ;
		star_id:_FillValue = -1s ;
		star_id:coordinates = "band_id band_wavelength_star_look t_star_look" ;
	int channel_integration_time ;
		channel_integration_time:long_name = "Channel-dependent Channel Integration Time, as defined in the VNIR or IR Channel Configuration Table Telemetry" ;
		channel_integration_time:_FillValue = -1 ;
		channel_integration_time:units = "count" ;
	int channel_gain_field ;
		channel_gain_field:long_name = "Channel-dependent Gain Field, as defined in the VNIR or IR Channel Configuration Table Telemetry" ;
		channel_gain_field:_FillValue = -1 ;
		channel_gain_field:units = "1" ;

// global attributes:
		:naming_authority = "gov.nesdis.noaa" ;
		:Conventions = "CF-1.7" ;
		:standard_name_vocabulary = "CF Standard Name Table (v35, 20 July 2016)" ;
		:institution = "DOC/NOAA/NESDIS > U.S. Department of Commerce, National Oceanic and Atmospheric Administration, National Environmental Satellite, Data, and Information Services" ;
		:project = "GOES" ;
		:production_site = "WCDAS" ;
		:production_environment = "OE" ;
		:spatial_resolution = "1km at nadir" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:orbital_slot = "GOES-East" ;
		:platform_ID = "G16" ;
		:instrument_type = "GOES-R Series Advanced Baseline Imager (ABI)" ;
		:scene_id = "Full Disk" ;
		:instrument_ID = "FM1" ;
		:title = "ABI L1b Radiances" ;
		:summary = "Single reflective band ABI L1b Radiance Products are digital maps of outgoing radiance values at the top of the atmosphere for visible and near-IR bands." ;
		:keywords = "SPECTRAL/ENGINEERING > VISIBLE WAVELENGTHS > VISIBLE RADIANCE" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Earth Science Keywords, Version 7.0.0.0.0" ;
		:iso_series_metadata_id = "a70be540-c38b-11e0-962b-0800200c9a66" ;
		:license = "Unclassified data.  Access is restricted to approved users only." ;
		:processing_level = "National Aeronautics and Space Administration (NASA) L1b" ;
		:cdm_data_type = "Image" ;
		:dataset_name = "OR_ABI-L1b-RadF-M6C01_G16_s20220011800205_e20220011809513_c20220011809562.nc" ;
		:production_data_source = "Realtime" ;
		:timeline_id = "ABI Mode 6" ;
		:date_created = "2022-01-01T18:09:56.2Z" ;
		:time_coverage_start = "2022-01-01T18:00:20.5Z" ;
		:time_coverage_end = "2022-01-01T18:09:51.3Z" ;
		:LUT_Filenames = "SpaceLookParams(FM1A_CDRL79RevP_PR_09_00_02)-637827000.0.h5 QTableBand01(FM1A_CDRL79RevH_DO_07_00_00)-582860861.0.h5 CalTargetTimeIntervals(FM1A_CDRL79RevP_DO_08_00_01)-611906620.0.h5 BandSaturationLimits(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.h5 SolarSpaceLookParams(FM1A_CDRL79RevH_DO_09_00_00)-600765435.0.h5 DeadRowListParams(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.h5 Mirror_Record(FM1A_CDRL79RevG_DO_07_00_00)-582860861.0.h5 KalmanAstroConsts(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.xml KalmanFilterControls(FM1A_PR_09_08_02)-677650371.0.xml KalmanMeasMaxSensibles(FMAA_INT_ONLY_DO_09_01_00)-652936814.0.xml KalmanPreprocessorControls(FM1A_CDRL79RevJ_PR_09_06_02)-657795700.0.xml KalmanReferenceData(FM1A_CDRL79RevH_DO_08_00_00)-888.0.xml KalmanStarCatalogs(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.xml ABI_NavigationRDP_Band01(FM1A_CDRL79RevJ_DO_07_00_00)-582860861.0.xml ABI_NavigationParameters_Band01(FM1A_CDRL79RevH_DO_07_00_00)-582860861.0.xml ABI_ResamplingImplementation_Band01(FM1A_CDRL79RevH_DO_07_02_00)-602129336.0.xml ABI_ResamplingParameters_Band01(FM1A_CDRL79RevJ_DO_07_00_00)-582860861.0.xml StarLookParams(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.h5 StarDetectionParams(FM1A_CDRL79RevJ_DO_07_00_00)-582860861.0.xml ResamplingScaledConversion(FMAA_INT_ONLY_DO_08_00_00)-1111.0.xml BlockReleaseRegions(FMAA_INT_ONLY_DO_08_00_00)-2222.0.csv VNIR_RetrievalParameters(FM1A_CDRL79RevH_DO_08_00_00)-600000000.0.h5 SCT_Record(FM1A_CDRL79RevM_DO_09_00_00)-600765435.0.h5 ICM_ConversionConsts(FM1A_CDRL43-18_DO_09_01_00)-652936750.0.h5 ICM_SensorCoefficients(FM1A_TMABI_18_159_TMABI_18_533_DO_09_05_00)-676949608.0.h5" ;
		:id = "75de858d-c386-4159-a95e-bce8a0d3d61e" ;
}
