[0] /.zgroup : (50) |{
"foo": 42,
"bar": "apples",
"baz": [1, 2, 3, 4]}|
[1] /meta1/.zarray : (34) |{
"shape": [1,2,3],
"dtype": "<1"}|
