netcdf ref_tst_nul3 {
dimensions:
	n = 8 ;
variables:
	char cdata(n) ;
	char c;

// global attributes:
		:global = "x\000y" ;
data:

 cdata = "abc\000def" ;

 c = "";
}
