netcdf appel {
types:
  int(*) vlen_int ;
  compound singleCompoundType {
    vlen_int vlenIntVector(2) ;
  }; // singleCompoundType
  compound pfCoilType {
    vlen_int name ;
  }; // pfCoilType
  pfCoilType(*) vlen_t ;
  vlen_int(*) vlen_int2 ;
  compound singleCompoundType2 {
    vlen_int2 vlenIntVector ;
  }; // singleCompoundType2
dimensions:
	vlenDim = 2 ;
variables:
	vlen_int vdata ;
	singleCompoundType singleCompound ;
	vlen_t pfCircuits ;
	singleCompoundType2 singleCompound2 ;
	vlen_int vlenIntVector(vlenDim) ;
data:

 vdata = {1, 2, 3} ;

 singleCompound = {{{11}, {12}}} ;

 pfCircuits = {{{1, 2, 3}}, {{2}}, {{3}}, {{4}}} ;

 singleCompound2 = {{{11}, {12}}} ;

 vlenIntVector = {1, 2, 3}, {1, 2, 3} ;
}
