[0] /.zgroup : (0) ||
[1] /meta1/.zarray : (50) |{
"foo": 42,
"bar": "apples",
"baz": [1, 2, 3, 4]}|
[2] /meta2/.zarray : (64) |{
"foo": 42,
"bar": "apples",
"baz": [1, 2, 3, 4],
"extra": 137}|
