netcdf testmeta {

group: _nczarr {

  // group attributes:
  		:data = "{\"zarr_format\": 2,\"nczarr_version\": \"1.0.0\"}" ;
  } // group _nczarr

group: _zgroup {

  // group attributes:
  		:data = "{\"zarr_format\": 2}" ;
  } // group _zgroup

group: _nczgroup {

  // group attributes:
  		:data = "{\"dimensions\": {},\"arrays\": [\"var1\"],\"groups\": []}" ;
  } // group _nczgroup

group: _nczattr {

  // group attributes:
  		:data = "{\"types\": {\"_NCProperties\": \"2\"}}" ;
  } // group _nczattr

group: _zattrs {

  // group attributes:
  		:data = "{\"_NCProperties\": \"version=\"}" ;
  } // group _zattrs

group: var1 {

  group: _zarray {

    // group attributes:
    		:data = "{\"zarr_format\": 2,\"shape\": [],\"dtype\": \"<i4\",\"chunks\": [],\"fill_value\": -2147483647,\"order\": \"C\",\"compressor\": null,\"filters\": null}" ;
    } // group _zarray

  group: _nczvar {

    // group attributes:
    		:data = "{\"dimension_references\": [],\"contiguous\": true}" ;
    } // group _nczvar
  } // group var1
}
