netcdf test_test {

types:
  byte enum enum_t {c1=1, c2=2, c3=3};

variables:
  enum_t v1;

data:
  v1 = c1;
}
