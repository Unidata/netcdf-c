netcdf tst_mud4 {
dimensions:
	F0 = 1 ;
	F1 = 2 ;
	F2 = 3 ;
	F3 = 5 ;
	U0 = UNLIMITED ; // (1 currently)
	U1 = UNLIMITED ; // (2 currently)
	U2 = UNLIMITED ; // (3 currently)
	U3 = UNLIMITED ; // (5 currently)
variables:
	int ff(F1, F2) ;
		ff:_FillValue = -2147483647 ;
	int uf(U1, F2) ;
		uf:_FillValue = -2147483647 ;
	int fu(F1, U2) ;
		fu:_FillValue = -2147483647 ;
	int uu(U1, U2) ;
		uu:_FillValue = -2147483647 ;
	int ufff(U0, F1, F2, F3) ;
		ufff:_FillValue = -2147483647 ;
	int uffu(U0, F1, F2, U3) ;
		uffu:_FillValue = -2147483647 ;
	int ufuf(U0, F1, U2, F3) ;
		ufuf:_FillValue = -2147483647 ;
	int ufuu(U0, F1, U2, U3) ;
		ufuu:_FillValue = -2147483647 ;
	int uuff(U0, U1, F2, F3) ;
		uuff:_FillValue = -2147483647 ;
	int uufu(U0, U1, F2, U3) ;
		uufu:_FillValue = -2147483647 ;
	int uuuf(U0, U1, U2, F3) ;
		uuuf:_FillValue = -2147483647 ;
	int uuuu(U0, U1, U2, U3) ;
		uuuu:_FillValue = -2147483647 ;
	int ffff(F0, F1, F2, F3) ;
		ffff:_FillValue = -2147483647 ;
data:

 ff =
  1, 2, 3,
  4, 5, 6 ;

 uf =
  1, 2, 3,
  4, 5, 6 ;

 fu =
  {1, 2, 3},
  {4, 5, 6} ;

 uu =
  {1, 2, 3},
  {4, 5, 6} ;

 ufff =
  1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30 ;

 uffu =
  {1, 2, 3, 4, 5},
  {6, 7, 8, 9, 10},
  {11, 12, 13, 14, 15},
  {16, 17, 18, 19, 20},
  {21, 22, 23, 24, 25},
  {26, 27, 28, 29, 30} ;

 ufuf =
  {1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15},
  {16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30} ;

 ufuu =
  {{1, 2, 3, 4, 5},
  {6, 7, 8, 9, 10},
  {11, 12, 13, 14, 15}},
  {{16, 17, 18, 19, 20},
  {21, 22, 23, 24, 25},
  {26, 27, 28, 29, 30}} ;

 uuff =
  {1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30} ;

 uufu =
  {{1, 2, 3, 4, 5},
  {6, 7, 8, 9, 10},
  {11, 12, 13, 14, 15},
  {16, 17, 18, 19, 20},
  {21, 22, 23, 24, 25},
  {26, 27, 28, 29, 30}} ;

 uuuf =
  {{1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15},
  {16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30}} ;

 uuuu =
  {{{1, 2, 3, 4, 5},
  {6, 7, 8, 9, 10},
  {11, 12, 13, 14, 15}},
  {{16, 17, 18, 19, 20},
  {21, 22, 23, 24, 25},
  {26, 27, 28, 29, 30}}} ;

 ffff =
  1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30 ;
}
