[1] /.nczarr : (0) ||
