netcdf n3time {
dimensions:
	Mode = 10 ;
	NameLength = 32 ;
	Heights = 69 ;
	SpectraPoints = 256 ;
	TimeSeriesPoints = 12288 ;
	Beams = 5 ;
	Time = UNLIMITED ; // (10 currently)
variables:
	char DwellModeName(Mode, NameLength) ;
		DwellModeName:long_name = "Name of the dwell mode" ;
	float ClutterHeight(Mode) ;
		ClutterHeight:long_name = "Maximum height of clutter removal" ;
		ClutterHeight:units = "meters" ;
	short ClutterRemovedGates(Mode) ;
		ClutterRemovedGates:long_name = "Number of gates removed by clutter algorithm" ;
		ClutterRemovedGates:units = "count" ;
	short CodeBits(Mode) ;
		CodeBits:long_name = "Number of code bits" ;
		CodeBits:units = "count" ;
	short CoherentIntegrations(Mode) ;
		CoherentIntegrations:long_name = "Number of coherent integrations" ;
		CoherentIntegrations:units = "count" ;
	short ConcatenatedTimeSeries(Mode) ;
		ConcatenatedTimeSeries:long_name = "Concatenated time series" ;
		ConcatenatedTimeSeries:units = "0 = off, 1 = on" ;
	short DcFilterOn(Mode) ;
		DcFilterOn:long_name = "Spectral filtering of DC" ;
		DcFilterOn:units = "0 = off, 1 = on" ;
	short DcOmittedPoints(Mode) ;
		DcOmittedPoints:long_name = "Number of points omitted around DC" ;
		DcOmittedPoints:units = "count" ;
	short DwellTimeConvention(Mode) ;
		DwellTimeConvention:long_name = "Dwell time convention" ;
		DwellTimeConvention:units = "0=begin,1=mid,2=end" ;
	int FirstGate(Mode) ;
		FirstGate:long_name = "Delay period to first range gate" ;
		FirstGate:units = "ns" ;
	float FirstHeight(Mode) ;
		FirstHeight:long_name = "Height of first range gat" ;
		FirstHeight:units = "meters" ;
	short Flip(Mode) ;
		Flip:long_name = "Phase flip DC removal" ;
		Flip:units = "0 = off, 1 = on" ;
	short Gates(Mode) ;
		Gates:long_name = "Number of range gates" ;
		Gates:units = "count" ;
	int GateSpacing(Mode) ;
		GateSpacing:long_name = "Height spacing of range gates" ;
		GateSpacing:units = "ns" ;
	float HeightSpacing(Mode) ;
		HeightSpacing:long_name = "Gate spacing" ;
		HeightSpacing:units = "meters" ;
	int InterPulsePeriod(Mode) ;
		InterPulsePeriod:long_name = "Inter-pulse period" ;
		InterPulsePeriod:units = "ns" ;
	float NyquistFrequency(Mode) ;
		NyquistFrequency:long_name = "Nyquist frequency" ;
		NyquistFrequency:units = "meters/second" ;
	short Overlap(Mode) ;
		Overlap:long_name = "Spectra" ;
		Overlap:units = "0 = off, 1 = on" ;
	int PreBlank(Mode) ;
		PreBlank:long_name = "Blank period before the transmit pulse" ;
		PreBlank:units = "ns" ;
	int PreTR(Mode) ;
		PreTR:long_name = "TR period before the transmit pulse" ;
		PreTR:units = "ns" ;
	int PostBlank(Mode) ;
		PostBlank:long_name = "Blank period after the transmit pulse" ;
		PostBlank:units = "ns" ;
	int PostTR(Mode) ;
		PostTR:long_name = "TR period after the transmit pulse" ;
		PostTR:units = "ns" ;
	int RassBeginPoint(Mode) ;
		RassBeginPoint:long_name = "First RASS spectral point" ;
		RassBeginPoint:units = "count" ;
	short RassHighFrequency(Mode) ;
		RassHighFrequency:long_name = "Upper frequency of RASS audio source" ;
		RassHighFrequency:units = "Hz" ;
	short RassLowFrequency(Mode) ;
		RassLowFrequency:long_name = "Lower frequency of RASS audio source" ;
		RassLowFrequency:units = "Hz" ;
	short RassOn(Mode) ;
		RassOn:long_name = "RASS On" ;
		RassOn:units = "0 = off, 1 = on" ;
	int RassPoints(Mode) ;
		RassPoints:long_name = "Number of RASS spectral points" ;
		RassPoints:units = "count" ;
	short RassStep(Mode) ;
		RassStep:long_name = "Step frequency of RASS audio source" ;
		RassStep:units = "Hz" ;
	short RassStepPeriod(Mode) ;
		RassStepPeriod:long_name = "Step period of RASS audio source" ;
		RassStepPeriod:units = "ns" ;
	short RassSweep(Mode) ;
		RassSweep:long_name = "RASS sweep type" ;
		RassSweep:units = "0 = random, 1 = sweep" ;
	int ReceiverDelay(Mode) ;
		ReceiverDelay:long_name = "Receiver delay period" ;
		ReceiverDelay:units = "ns" ;
	short ReceiverMode(Mode) ;
		ReceiverMode:long_name = "Receiver mode" ;
		ReceiverMode:units = "0 = multiple antennas, 1 = dual polarization" ;
	short Receivers(Mode) ;
		Receivers:long_name = "Number of receiver" ;
		Receivers:units = "count" ;
	short SpectralAverages(Mode) ;
		SpectralAverages:long_name = "Number of spectral averages" ;
		SpectralAverages:units = "count" ;
	short SpectralAverageType(Mode) ;
		SpectralAverageType:long_name = "Spectral average type" ;
		SpectralAverageType:units = "0 = mean, 1 = ICRA" ;
	int SpectralPoints(Mode) ;
		SpectralPoints:long_name = "Number of points in FFT" ;
		SpectralPoints:units = "count" ;
	int TxPulseWidth(Mode) ;
		TxPulseWidth:long_name = "Transmit pulse duration" ;
		TxPulseWidth:units = "ns" ;
	short VerticalCorrectHw(Mode) ;
		VerticalCorrectHw:long_name = "Vertical correction implemented in hardware" ;
		VerticalCorrectHw:units = "0 = off, 1 = on" ;
	float VerticalCorrectHwAngle(Mode) ;
		VerticalCorrectHwAngle:long_name = "Elevation angle used in hardware vertical correction" ;
		VerticalCorrectHwAngle:units = "degrees" ;
	int WindBeginPoint(Mode) ;
		WindBeginPoint:long_name = "First wind spectral point" ;
		WindBeginPoint:units = "count" ;
	int WindPoints(Mode) ;
		WindPoints:long_name = "Number Of wind spectral points" ;
		WindPoints:units = "count" ;
	short WindowingType(Mode) ;
		WindowingType:long_name = "Spectral window type" ;
		WindowingType:units = "0 = no window, 1 = Hann" ;
	short ModeNumber(Time) ;
		ModeNumber:long_name = "NetCDF index for dwell mode parameter sets" ;
		ModeNumber:units = "count" ;
	float Latitude(Time) ;
		Latitude:long_name = "Latitude of radar" ;
		Latitude:units = "degrees north" ;
	float Longitude(Time) ;
		Longitude:long_name = "Longitude of radar" ;
		Longitude:units = "degrees east" ;
	int Altitude(Time) ;
		Altitude:long_name = "Altitude of radar" ;
		Altitude:units = "meters above sea level" ;
	float Azimuth(Time) ;
		Azimuth:long_name = "Azimuth angle of the beam of the array" ;
		Azimuth:units = "degrees" ;
	float Elevation(Time) ;
		Elevation:long_name = "Elevation angle of the beam of the array" ;
		Elevation:units = "degrees" ;
	int DirectionCode(Time) ;
		DirectionCode:long_name = "Direction code of" ;
		DirectionCode:units = "count" ;
	char BeamDirection(Time, NameLength) ;
		BeamDirection:long_name = "Direction of beam" ;
	int Timestamp(Time) ;
		Timestamp:long_name = "Time in Unix Epoch" ;
		Timestamp:units = "seconds since 1970-1-1 0:00:00 0:00" ;
	int TimestampMilliseconds(Time) ;
		TimestampMilliseconds:long_name = "Milliseconds offset from timestamp" ;
		TimestampMilliseconds:units = "milliseconds" ;
	float MeanDopplerVelocity(Time, Heights) ;
		MeanDopplerVelocity:long_name = "Mean Doppler velocity" ;
		MeanDopplerVelocity:units = "meters/sec" ;
		MeanDopplerVelocity:missing_value = "9.9692099683868690e+36" ;
	float SNR(Time, Heights) ;
		SNR:long_name = "Signal to noise ratio" ;
		SNR:units = "dB" ;
		SNR:missing_value = "9.9692099683868690e+36" ;
	float Power(Time, Heights) ;
		Power:long_name = "Power" ;
		Power:units = "dB" ;
		Power:missing_value = "9.9692099683868690e+36" ;
	float SpectralWidth(Time, Heights) ;
		SpectralWidth:long_name = "Spectral width" ;
		SpectralWidth:units = "meters/sec" ;
		SpectralWidth:missing_value = "9.9692099683868690e+36" ;
	float NoiseLevel(Time, Heights) ;
		NoiseLevel:long_name = "Mean noise level" ;
		NoiseLevel:units = "dB" ;
		NoiseLevel:missing_value = "9.9692099683868690e+36" ;

// global attributes:
		:StationID = "BOU_DEMO_LAP161" ;
		:StationName = "LAP161 Demonstration" ;
		:RadarID = 2009 ;
		:WMOStationNumber = -1 ;
		:Location = "Louisville, Colorado" ;
		:AlignmentDeg = 0.f ;
		:LapxmVersion = "2.5.0.0" ;
		:ConfigFile = "NetCDF4 10.cfg" ;
		:DataTypes = "Moments," ;
		:TimeOfFirstRecord = "07-Apr-2009,17:43:17 GMT" ;
		:MinutesToUTC = 360s ;
data:

 DwellModeName =
  "WA",
  "WB",
  "WC",
  "WD",
  "WE",
  "WF",
  "WG",
  "WH",
  "WI",
  "WJ" ;

 ClutterHeight = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 ClutterRemovedGates = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 CodeBits = 1, 4, 1, 4, 1, 4, 1, 4, 1, 4 ;

 CoherentIntegrations = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

 ConcatenatedTimeSeries = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DcFilterOn = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 DcOmittedPoints = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 DwellTimeConvention = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FirstGate = 4083, 23000, 4083, 23000, 4083, 23000, 4083, 23000, 4083, 23000 ;

 FirstHeight = 188.6541, 2344.907, 188.6541, 2344.907, 188.6541, 2344.907, 
    188.6541, 2344.907, 188.6541, 2344.907 ;

 Flip = 1, 0, 1, 0, 1, 0, 1, 0, 1, 0 ;

 Gates = 60, 61, 62, 63, 64, 65, 66, 67, 68, 69 ;

 GateSpacing = 667, 1333, 667, 1333, 667, 1333, 667, 1333, 667, 1333 ;

 HeightSpacing = 96.49825, 192.9965, 96.49825, 192.9965, 96.49825, 192.9965, 
    96.49825, 192.9965, 96.49825, 192.9965 ;

 InterPulsePeriod = 93000, 151000, 93000, 151000, 93000, 151000, 93000, 
    151000, 93000, 151000 ;

 NyquistFrequency = 897.4543, 552.7368, 897.4543, 552.7368, 897.4543, 
    552.7368, 897.4543, 552.7368, 897.4543, 552.7368 ;

 Overlap = 1, 0, 1, 0, 1, 0, 1, 0, 1, 0 ;

 PreBlank = 3000, 3000, 3000, 3000, 3000, 3000, 3000, 3000, 3000, 3000 ;

 PreTR = 1500, 1500, 1500, 1500, 1500, 1500, 1500, 1500, 1500, 1500 ;

 PostBlank = 1500, 2500, 1500, 2500, 1500, 2500, 1500, 2500, 1500, 2500 ;

 PostTR = 396, 396, 396, 396, 396, 396, 396, 396, 396, 396 ;

 RassBeginPoint = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 RassHighFrequency = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 RassLowFrequency = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 RassOn = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RassPoints = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RassStep = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 RassStepPeriod = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 RassSweep = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1 ;

 ReceiverDelay = 2780, 6800, 2780, 6800, 2780, 6800, 2780, 6800, 2780, 6800 ;

 ReceiverMode = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Receivers = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 SpectralAverages = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 ;

 SpectralAverageType = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 SpectralPoints = 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024 ;

 TxPulseWidth = 1000, 5333, 1000, 5333, 1000, 5333, 1000, 5333, 1000, 5333 ;

 VerticalCorrectHw = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 VerticalCorrectHwAngle = 75, 75, 75, 75, 75, 75, 75, 75, 75, 75 ;

 WindBeginPoint = 384, 384, 384, 384, 384, 384, 384, 384, 384, 384 ;

 WindPoints = 256, 256, 256, 256, 256, 256, 256, 256, 256, 256 ;

 WindowingType = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ModeNumber = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 Latitude = 39.97, 39.97, 39.97, 39.97, 39.97, 39.97, 39.97, 39.97, 39.97, 
    39.97 ;

 Longitude = -105.12, -105.12, -105.12, -105.12, -105.12, -105.12, -105.12, 
    -105.12, -105.12, -105.12 ;

 Altitude = 1634, 1634, 1634, 1634, 1634, 1634, 1634, 1634, 1634, 1634 ;

 Azimuth = 90, 0, 270, 270, 0, 90, 90, 0, 270, 90 ;

 Elevation = 90, 75, 75, 75, 75, 90, 90, 75, 75, 90 ;

 DirectionCode = 1, 2, 3, 3, 2, 1, 1, 2, 3, 1 ;

 BeamDirection =
  "Vertical",
  "North",
  "West",
  "West",
  "North",
  "Vertical",
  "Vertical",
  "North",
  "West",
  "Vertical" ;

 Timestamp = 1239126197, 1239126199, 1239126200, 1239126202, 1239126203, 
    1239126205, 1239126207, 1239126208, 1239126210, 1239126212 ;

 TimestampMilliseconds = 466, 138, 779, 341, 982, 545, 201, 857, 404, 14 ;

 MeanDopplerVelocity =
  43.82101, 58.27499, 72.74288, 87.21077, 101.6647, 116.1187, 130.5866, 
    145.0545, 159.5085, 173.9625, 188.4304, 202.8982, 217.3522, 219.1318, 
    215.5473, 211.3465, 197.2325, 204.179, 196.8286, 188.8497, 178.6756, 
    203.4626, 150.1544, 146.7364, 161.4521, 59.54426, 80.96873, 95.59282, 
    184.9923, -0.00545623, 0.01037753, 52.64631, 145.692, 0.01144738, 
    -0.004172411, 0.01048452, 115.5366, 0.01230326, -0.06140933, -0.01406851, 
    171.7784, -0.03637486, -0.005349245, 0.02289477, -218.4591, -0.03016974, 
    0.03594692, 0.007274973, -159.5085, -0.0311326, -0.03546549, 0.004065426, 
    -99.91191, -0.01144738, 0.0148709, -0.01144738, -42.06817, -0.01299866, 
    -0.004493366, 0.007916883, _, _, _, _, _, _, _, _, _,
  26.9891, 35.62561, 44.26212, 52.89864, 61.53514, 70.17166, 78.80817, 
    87.44468, 96.08119, 104.7177, 113.3542, 121.9907, 130.6272, 135.1799, 
    130.9728, 126.9807, 123.3603, 119.8915, 116.8655, 114.0557, 111.0854, 
    108.4877, 106.6398, 104.6201, 102.2249, 101.6468, 99.74647, 99.24543, 
    96.17548, 94.32571, 115.2055, 111.2, 92.35497, 89.6981, 89.6162, 53.9782, 
    62.61471, 123.103, 77.72861, 119.1437, 119.1735, 106.9307, 121.8901, 
    121.9907, 130.6035, -136.0251, -129.5477, -119.8316, -111.1951, -101.479, 
    -95.00163, -85.28555, -77.72861, 134.962, -59.38808, 88.52425, -43.18256, 
    -32.38692, -24.82997, -17.27302, -6.477384, _, _, _, _, _, _, _, _,
  43.82101, 57.84374, 71.86646, 85.88918, 99.91191, 113.9346, 127.9574, 
    141.9801, 156.0028, 170.0255, 184.0482, 198.071, 212.0937, 219.4856, 
    212.655, 206.1729, 200.2946, 194.6629, 189.7493, 185.1881, 180.3644, 
    176.1251, 173.1675, 169.8671, 165.9478, 165.0351, 161.9574, 161.1433, 
    156.1496, 153.3434, 187.0545, 180.5443, 149.9528, 145.692, 145.453, 
    87.64203, 101.6647, 199.8747, 126.2045, 184.0934, 193.4987, 173.6212, 
    197.8694, 198.071, 212.0562, -220.8579, -210.3409, -194.5653, -180.5426, 
    -164.767, -154.25, -138.4744, -126.2045, 219.1332, -96.42575, 143.7329, 
    -70.11362, -52.58522, 15.77556, -28.04545, -10.51704, 2.203247, _, _, _, 
    _, _, _, _,
  26.9891, 35.36, 43.72234, 52.08896, 60.45558, 68.8222, 77.18883, 85.55544, 
    93.92207, 102.2887, 110.6553, 119.0219, 127.3885, 135.655, 134.8579, 
    133.313, 125.0804, 127.5444, 125.3105, 128.8786, 113.6978, 112.6653, 
    104.8687, 0.01917438, 104.9029, 86.49361, 0.01080618, 0.01844958, 
    97.27106, 55.63919, 0.000922479, 0.0007248049, 111.2, 0.003755807, 
    0.0003953481, -0.004085264, 52.89864, -0.006391461, 6.036703, 
    0.003294568, 86.36512, 0.00342635, 0.004678286, 0.004217047, 119.3348, 
    0.01186044, 0.05277898, -0.0144961, -124.1499, 0.006062005, 0.001581392, 
    0.001054262, -91.76294, -0.0263236, 0.01930617, 0.001383718, 80.91775, 
    -0.01186044, -0.006424407, 0, -24.82997, 0.03729451, 0.005600765, _, _, 
    _, _, _, _,
  43.82101, 57.41248, 70.99004, 84.57455, 98.15907, 111.7436, 125.3281, 
    138.9057, 152.4971, 166.0886, 179.6662, 193.2507, 206.8352, 220.257, 
    218.9629, 216.4544, 203.0871, 207.0907, 203.4669, 209.2478, 184.6155, 
    182.8169, 170.2026, 0.02075507, 170.3237, 140.3428, 0.02214587, 
    0.01636869, 157.9315, 90.85446, -0.02567638, 0.02310874, 180.5443, 
    52.64631, -0.0009093716, -0.00962864, 85.88918, -0.01358708, 
    -0.006633063, 0.005777184, 140.2272, 0.01947125, -0.02235984, 
    -0.004065426, 193.7595, 0.02043412, 0.06857732, -0.01390804, -201.5767, 
    -0.006151631, -0.008772762, -0.00460035, -148.9914, -0.02524843, 
    0.03252341, 0.005563214, 131.3866, -0.01283819, -0.02749512, 0.00524226, 
    -40.31533, 0.09757023, 0.002781607, 0.06847033, _, _, _, _, _,
  26.9891, 35.08583, 43.18256, 51.27929, 59.37602, 67.47275, 75.56948, 
    83.66621, 91.76294, 99.85966, 107.9564, 116.0531, 124.1499, 132.2465, 
    134.6545, 133.9732, 126.9807, 129.3814, 120.3224, 124.0806, 114.4163, 
    115.755, 110.035, 124.8917, 104.5875, 0.0001317827, 101.4128, 
    0.004217047, 116.6242, 46.55132, 96.53848, 0.000922479, 115.2055, 
    0.007841071, 119.5976, 0.01001549, 87.07576, 0.003953482, 118.6575, 
    -0.02095345, 74.6209, 0.01304649, 92.19202, -0.007412778, 105.7973, 
    0.00144961, 122.7255, 0.01396897, -136.0251, -0.001713175, -121.7413, 
    0.009751921, -104.7177, -0.004184101, -89.60381, -0.01887787, -72.33079, 
    0.02299608, 82.0547, -0.006062005, -39.56908, -0.03765691, -24.82997, 
    0.01205812, -6.477384, _, _, _, _,
  43.82101, 56.96732, 70.11362, 83.25993, 96.40623, 109.5525, 122.6988, 
    135.8451, 148.9914, 162.1377, 175.2841, 188.4304, 201.5767, 214.723, 
    218.6326, 216.853, 206.1729, 210.0725, 195.3589, 201.4607, 185.7733, 
    187.9821, 178.6756, 166.8432, 169.8126, 137.9689, 164.6606, 105.1839, 
    189.3544, 75.59274, 156.7598, -0.02567638, 187.0545, 0.01037753, 
    194.1849, 0.02000618, 141.3645, 0.0170106, 192.6556, -0.004065426, 
    121.1707, 0.01358708, 149.6873, -0.02203889, 171.7784, 3.120749, 
    199.2624, 0.02161095, -220.8579, 0.006954018, -197.6698, 0.008986731, 
    -170.0255, -0.008665777, -145.4858, -0.03546549, -117.4403, 0.002781607, 
    133.2279, -0.003851456, -64.24641, -0.03551899, -40.31533, 0.01315914, 
    -10.51704, 0.01925728, _, _, _,
  26.9891, 34.81166, 42.64278, 50.4739, 58.29646, 66.12329, 73.95013, 
    81.78126, 89.60381, 97.43065, 105.2575, 113.0843, 120.9112, 128.7337, 
    136.0251, 134.7499, 128.9336, 132.049, 128.4584, 125.3424, 116.1737, 
    127.9053, 114.3732, 109.8473, 106.9696, 0.02194182, 83.74001, 84.40551, 
    101.0611, 0.01462788, 46.55132, 55.63919, 94.32571, -0.00342635, 
    0.009158898, 0.02892631, 92.85463, 0.01008138, -0.001317827, 
    -0.004282938, 64.77384, -0.04958325, -0.003228677, -0.008829442, 
    96.08119, -0.01535269, 0.0002635654, -0.006193787, 125.2294, 
    0.0003953481, -0.0144961, -0.01080618, -119.8316, 0.00632557, 
    -0.0002635654, -0.009718975, -88.52425, -0.01759299, -0.0350542, 
    0.03571311, 82.0547, -0.0003294568, -0.006424407, 0.02503872, -24.82997, 
    -0.004777123, 0.01429842, _, _,
  43.82101, 56.52215, 69.2372, 81.95225, 94.65339, 107.3615, 120.0696, 
    132.7846, 145.4858, 158.1939, 170.9019, 183.617, 196.3181, 209.0262, 
    220.7865, 218.7875, 209.3436, 214.4024, 208.5739, 203.5288, 188.626, 
    207.6793, 185.6689, 178.3787, 173.6824, 0.02931386, 135.8394, 136.9278, 
    164.0877, 0.01112643, 75.59274, 90.85446, 153.3434, -0.00545623, 
    0.007809897, 55.23545, 150.7582, -0.003583994, -0.01027055, 1.123555, 
    105.1704, -0.07242877, -0.007061003, 0.01230326, 156.0028, -0.007167988, 
    -0.005723692, -0.02364366, 203.3295, -0.01305216, -0.01604773, 
    -0.003958441, -194.5653, -0.00545623, 0.002460652, -0.009682133, 
    -143.7329, -0.01829442, -0.04787574, 0.03091864, 133.2279, 0.003423517, 
    -0.02749512, 0.02139698, 15.77556, 0.002567637, -0.004493366, 
    -0.04290094, _,
  26.9891, 34.54605, 42.103, 49.65994, 57.21689, 64.77384, 72.33079, 
    79.88773, 87.44468, 95.00163, 102.5586, 110.1155, 117.6725, 125.2294, 
    132.7864, 134.6545, 130.9728, 127.4628, 124.1521, 120.9648, 118.1041, 
    115.1428, 113.0708, 110.91, 108.4877, 106.4837, 104.1555, 101.8097, 
    100.8984, 101.0611, 116.6242, 97.27106, 96.17548, 113.9356, 115.5939, 
    91.35184, 115.5704, 121.2415, 89.53384, 46.42125, 53.9782, 61.53514, 
    116.7609, 117.3785, 83.12643, 92.19202, 99.66483, 104.7177, 121.8901, 
    120.9127, 128.8421, 134.9553, -131.7068, -124.1499, -117.6749, -110.1155, 
    -101.479, -96.08119, -88.52425, -80.9673, -72.33079, 73.41035, 80.91775, 
    88.52425, -43.18256, -34.54605, -25.90953, -18.35259, 126.309 ;

 SNR =
  73.58841, 93.69621, 90.72098, 93.79675, 73.58717, 95.86793, 69.22738, 
    97.28767, 73.58855, 104.8742, 101.2131, 103.8415, 76.61465, 66.12689, 
    51.4962, 36.75954, 17.05997, 43.50135, 30.1532, 21.94452, 9.951521, 
    14.91348, 23.56355, 15.50947, 7.67453, 23.93628, 20.8658, 13.8817, 
    -0.9981411, 13.75913, 4.403778, 13.87306, 4.132092, 15.36119, 7.184721, 
    2.787889, -10.59243, 21.66834, 10.08679, 5.269455, 32.43215, 17.2073, 
    12.63988, 6.887564, -6.582558, 16.96766, 26.28023, 9.15701, 36.32301, 
    15.8774, 26.87329, 11.01729, 37.94886, 15.25741, 17.61534, 12.92631, 
    39.29753, 15.34392, 25.4152, 13.9917, _, _, _, _, _, _, _, _, _,
  73.58841, 73.58746, 73.58705, 73.58668, 73.58678, 73.58697, 73.58717, 
    73.58771, 73.58835, 73.59007, 73.59528, 73.62238, 74.16414, 48.64612, 
    29.8039, 22.89784, 18.98489, 16.34667, 14.86743, 12.00373, 11.01264, 
    10.80821, 10.88415, 8.367054, 8.34943, 6.596746, 7.390163, 8.169736, 
    6.133302, 5.994343, -1.464175, -1.038825, 4.349963, 4.132089, 7.472332, 
    36.92896, 37.58608, -5.406899, 37.82778, -5.064863, -4.13306, -10.49347, 
    -6.046967, 39.84547, -9.53551, 39.95054, 41.36459, 41.64101, 41.68096, 
    43.30532, 43.02773, 43.00186, 43.56744, -14.29854, -4.054775, 45.51334, 
    45.49855, 44.71341, 45.27624, 45.88882, 45.7173, _, _, _, _, _, _, _, _,
  73.58841, 73.58746, 73.58705, 73.58668, 73.58678, 73.58697, 73.58717, 
    73.58771, 73.58835, 73.59007, 73.59528, 73.62238, 74.16414, 48.70594, 
    29.80793, 22.89856, 18.98499, 16.34634, 14.86528, 12.00291, 11.01402, 
    10.86728, 10.80384, 8.36587, 8.413319, 6.599803, 7.388638, 8.162623, 
    6.131635, 5.916479, -1.468702, -1.026616, 4.349304, 4.132092, 7.601118, 
    30.87293, 31.58507, -5.42053, 31.76128, -3.400933, -4.119135, -10.50972, 
    -6.032066, 33.80612, -9.534983, 33.95592, 35.35545, 35.59553, 35.65208, 
    37.26597, 36.98692, 36.97174, 37.48088, -14.21466, -4.023761, 39.31638, 
    39.43657, 38.71969, 39.49628, 39.84634, 39.6381, -6.649632, _, _, _, _, 
    _, _, _,
  73.58841, 93.79379, 70.49077, 70.08128, 73.58749, 70.86732, 92.79933, 
    69.41212, 73.58818, 70.1161, 100.177, 76.7963, 73.73407, 105.1306, 
    46.61544, 37.51689, 20.22619, 31.77058, 33.48387, 19.83179, 11.11092, 
    20.39005, 25.95015, 9.703699, 7.973179, 15.9146, 4.011011, 9.813317, 
    6.262893, 15.01544, 3.448323, 13.5082, -1.038825, 0.2162695, 6.663949, 
    15.66912, 37.45469, 2.843141, 27.06795, 17.38095, 37.83796, 4.466388, 
    11.20273, 17.26732, -13.22419, 7.085457, 13.27443, 16.65663, 41.33859, 
    8.584423, 15.61247, 16.61092, 44.10894, 10.7135, 16.98459, 15.80502, 
    -10.34921, 12.17531, 18.0534, 23.8835, 44.38044, 13.50732, 18.95304, _, 
    _, _, _, _, _,
  73.58841, 93.80248, 70.49077, 70.08122, 73.58749, 70.08294, 69.22593, 
    99.89193, 73.58818, 99.99556, 69.51709, 74.00417, 73.73407, 105.128, 
    46.76748, 37.86553, 20.22952, 31.55587, 32.87184, 20.04547, 11.06594, 
    20.36798, 24.15219, 9.441714, 7.973078, 15.71288, 4.4901, 9.579041, 
    6.256992, 13.65437, 2.987458, 13.24016, -1.026616, 13.87306, 6.196348, 
    15.6901, 31.40908, 2.556067, 9.031481, 16.171, 31.79919, 4.340066, 
    11.12574, 16.45714, -13.2033, 6.915856, 12.91424, 16.49553, 35.42617, 
    8.662317, 15.16352, 15.84185, 38.08039, 10.65039, 16.90429, 15.31706, 
    -10.39488, 12.41246, 18.0153, 14.36253, 38.35535, 18.85924, 18.78527, 
    14.75542, _, _, _, _, _,
  73.58841, 70.48653, 73.58761, 71.05208, 73.58694, 70.50192, 73.58733, 
    94.52415, 73.58789, 98.18135, 73.59155, 101.2159, 73.64521, 73.7626, 
    43.70144, 39.13026, 22.89784, 40.74371, 15.98459, 31.71367, 13.44021, 
    27.57239, 9.992734, 10.53715, 9.596519, 4.599466, 7.43125, 4.04748, 
    -0.1938949, 23.4408, 7.199106, 3.448323, -1.464175, 4.727225, -2.513843, 
    6.158762, 5.817806, 7.325817, -3.792603, 8.486688, -12.16173, 10.19361, 
    -12.83169, 10.87098, 38.43658, 12.2035, -10.9928, 13.38923, 39.95054, 
    14.55401, -6.104247, 14.99589, 42.15044, 15.99747, 42.91883, 27.76295, 
    43.4021, 17.7896, -6.730154, 18.48993, 5.23984, 18.3704, 44.38044, 
    18.28391, 45.7173, _, _, _, _,
  73.58841, 69.21068, 73.58761, 90.73901, 73.58694, 89.91195, 73.58733, 
    94.51604, 73.58789, 71.13646, 73.59155, 101.2131, 73.64521, 104.1776, 
    43.69957, 56.47713, 22.89856, 39.59184, 15.98874, 31.30631, 13.43907, 
    26.83986, 9.951521, 24.26562, 9.598264, 22.50379, 7.431938, 23.39528, 
    -0.1822964, 22.55742, 7.195879, 2.987458, -1.468702, 4.403778, -2.492411, 
    6.103886, 5.832101, 7.301615, -3.748032, 8.40478, -12.12319, 9.644305, 
    -12.84323, 10.67416, 32.43215, 26.07437, -11.02513, 13.0515, 33.95592, 
    14.36501, -6.134531, 15.09341, 36.13064, 16.1999, 36.79631, 26.87329, 
    37.40169, 26.11369, -6.678365, 17.96864, 5.051213, 18.35721, 38.35535, 
    18.35196, 39.6381, 19.41827, _, _, _,
  73.58841, 93.68493, 90.74884, 93.76166, 73.58714, 69.40633, 91.86413, 
    95.4968, 73.58786, 74.79911, 99.27956, 71.16159, 73.6159, 109.6338, 
    101.7956, 44.00277, 25.45438, 31.67448, 37.99788, 28.09372, 14.36661, 
    21.31573, 27.47247, 18.70392, 9.355213, 10.41595, 23.91235, 15.89867, 
    7.307194, 9.635264, 23.4408, 15.01544, 5.994343, 13.58617, 4.761446, 
    0.259647, 7.136021, 15.70831, 7.009398, 2.587076, 37.26254, 16.5996, 
    10.05981, 4.115768, 38.8725, 17.66912, 11.83648, 6.675002, 39.62537, 
    17.01511, 14.25439, 7.884811, 41.04591, 16.02794, 16.12646, 10.01866, 
    43.23695, 16.88727, 17.54112, 11.28917, -6.730154, 16.15187, 18.0534, 
    12.52568, 45.27624, 15.80998, 27.28624, _, _,
  73.58841, 93.6959, 70.4901, 93.77921, 73.58714, 72.23392, 91.87521, 
    95.49976, 73.58786, 71.53458, 99.27006, 101.9114, 73.6159, 74.1722, 
    72.05188, 43.92168, 25.45418, 30.97463, 37.4131, 28.06639, 14.36451, 
    20.36998, 27.44926, 18.70047, 9.353999, 11.0501, 22.18199, 15.55906, 
    7.306041, 9.510633, 22.55742, 13.65437, 5.916479, 13.75913, 4.376264, 
    14.48896, 7.127583, 15.23868, 6.797114, 15.34295, 31.26233, 16.23901, 
    10.11602, 3.923566, 32.8423, 17.1556, 11.74255, 6.258971, 33.58575, 
    16.96808, 13.80846, 8.085489, 35.02168, 15.80869, 15.4772, 9.982072, 
    37.20572, 16.33719, 17.0949, 11.37243, -6.678365, 15.88378, 18.0153, 
    12.33571, 39.49628, 15.33787, 25.4152, 14.27914, _,
  73.58841, 73.58763, 73.58725, 73.58718, 73.58704, 73.58717, 73.58721, 
    73.58759, 73.58771, 73.58845, 73.58965, 73.59292, 73.60313, 73.66388, 
    76.59731, 43.70144, 29.8039, 23.45033, 20.19151, 17.23576, 15.16196, 
    13.92838, 12.46472, 10.49867, 10.80821, 10.00584, 8.869205, 9.5312, 
    7.55749, 7.307194, -0.1938949, 6.262893, 6.133302, -0.9981267, -1.845291, 
    6.443112, -2.423464, -3.727809, 5.515008, 36.55381, 36.92896, 38.48117, 
    -3.615067, -3.617845, 36.94485, -12.83169, -10.50944, 38.32426, 
    -6.046967, -9.067388, -10.46475, -12.71363, 40.53381, 41.30886, 
    -8.024484, 41.42351, 43.30532, 43.20938, 43.23695, 42.9604, 43.4021, 
    44.82168, -10.34921, 45.18643, 45.49855, 45.50547, 45.22829, 45.45814, 
    45.43151 ;

 Power =
  43.90087, 43.88691, 43.89695, 43.88691, 43.90087, 43.88691, 43.90087, 
    43.88691, 43.90087, 43.88691, 43.89695, 43.88691, 43.90087, -15.93773, 
    -32.08697, -44.46257, -67.41553, -58.63432, -58.42065, -63.25468, 
    -77.16756, -74.04691, -69.35247, -72.06198, -82.86562, -78.93454, 
    -74.84628, -76.98456, -88.66276, -81.61904, -78.6766, -79.6946, -90.3644, 
    -82.42516, -79.35938, -82.34039, -101.5875, -82.99782, -80.04523, 
    -82.97546, -60, -83.52543, -80.52922, -83.49931, -101.3476, -83.90852, 
    -80.80966, -83.79858, -60, -84.15321, -81.06235, -84.1443, -60, 
    -84.33395, -81.28017, -84.30485, -60, -84.33688, -81.31423, -84.32729, _, 
    _, _, _, _, _, _, _, _,
  37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 
    37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, -40.28799, 
    -59.44931, -66.86259, -71.58028, -75.04754, -77.79921, -80.11113, 
    -82.09177, -83.80496, -85.33065, -86.77075, -88.07394, -89.30414, 
    -90.33333, -91.45734, -92.44866, -93.28663, -95.75604, -96.41407, 
    -95.89081, -96.38251, -97.33186, -60, -60, -103.3708, -60, -103.8217, 
    -104.5011, -110.0028, -106.33, -60, -110.007, -60, -60, -60, -60, -60, 
    -60, -60, -60, -120.4209, -109.6009, -60, -60, -60, -60, -60, -60, _, _, 
    _, _, _, _, _, _,
  43.90087, 43.90087, 43.90087, 43.90087, 43.90087, 43.90087, 43.90087, 
    43.90087, 43.90087, 43.90087, 43.90087, 43.90087, 43.90087, -34.26738, 
    -53.42873, -60.842, -65.55968, -69.02695, -71.77861, -74.09055, 
    -76.07129, -77.78339, -79.31123, -80.75031, -82.05192, -83.28357, 
    -84.31215, -85.43674, -86.42853, -87.27147, -89.73518, -90.39216, 
    -89.86938, -90.3644, -91.30737, -60, -60, -97.35206, -60, -96.84581, 
    -98.47652, -103.9909, -100.2988, -60, -103.9945, -60, -60, -60, -60, -60, 
    -60, -60, -60, -114.3961, -103.58, -60, -60, -60, -60, -60, -60, 
    -105.3947, _, _, _, _, _, _, _,
  37.88027, 37.86631, 37.88027, 37.88027, 37.88027, 37.88027, 37.87635, 
    37.88027, 37.88027, 37.88027, 37.87635, 37.88027, 37.88027, 37.56898, 
    -23.13032, -42.89674, -69.42675, -56.93001, -59.83706, -69.02055, 
    -80.90386, -71.30692, -72.50005, -85.65956, -87.14916, -78.85011, 
    -83.21961, -86.83295, -91.61378, -83.18546, -84.286, -87.68689, 
    -96.41407, -87.67651, -84.99927, -88.38306, -60, -88.31313, -85.31577, 
    -88.98383, -60, -88.99476, -86.19093, -89.6356, -112.1057, -89.39773, 
    -86.85876, -89.80238, -60, -89.76597, -86.96648, -90.13199, -60, 
    -90.14912, -87.16719, -90.31497, -115.7018, -90.33238, -87.25071, 
    -90.31918, -60, -90.32315, -87.38263, _, _, _, _, _, _,
  43.90087, 43.88691, 43.90087, 43.90087, 43.90087, 43.90087, 43.90087, 
    43.88691, 43.90087, 43.88691, 43.90087, 43.90087, 43.90087, 43.58958, 
    -17.10974, -36.87602, -63.4061, -50.90934, -53.81697, -62.99924, 
    -74.88372, -65.28799, -66.47926, -79.65327, -81.12852, -72.83289, 
    -77.19288, -80.81558, -85.59406, -77.17548, -78.2986, -81.64375, 
    -90.39216, -79.6946, -78.9618, -82.42593, -60, -82.29951, -79.60437, 
    -83.00989, -60, -82.97363, -80.12223, -83.55121, -106.0882, -83.38353, 
    -80.70398, -83.76965, -60, -83.78663, -80.91585, -84.12537, -60, 
    -84.10089, -81.15941, -84.32137, -109.6845, -84.27251, -81.25626, 
    -84.39972, -60, -84.24529, -81.37827, -84.01674, _, _, _, _, _,
  37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 
    37.87635, 37.88027, 37.87635, 37.88027, 37.87635, 37.88027, 37.88021, 
    -44.91081, -32.97261, -66.86259, -51.57779, -74.65687, -61.48507, 
    -79.59769, -68.18655, -83.18733, -74.27858, -86.10505, -82.69753, 
    -88.52267, -83.26312, -91.94852, -81.1367, -92.40703, -84.286, -95.75604, 
    -84.68906, -98.45298, -85.00283, -97.01009, -85.28387, -101.0442, 
    -85.54379, -108.4798, -85.87328, -111.9621, -86.13396, -60, -86.38757, 
    -110.8921, -86.52097, -60, -86.74469, -107.5268, -86.96725, -60, 
    -87.03231, -60, -87.0542, -60, -87.26109, -112.6061, -87.29953, 
    -109.9844, -87.39404, -60, -87.34997, -60, _, _, _, _,
  43.90087, 43.90087, 43.90087, 43.89695, 43.90087, 43.89695, 43.90087, 
    43.89695, 43.90087, 43.90087, 43.90087, 43.89695, 43.90087, 43.89695, 
    -38.89021, -26.84269, -60.842, -45.55724, -68.63626, -55.46424, 
    -73.57706, -62.16637, -77.16756, -67.04925, -80.08465, -70.65709, 
    -82.50203, -73.28304, -85.92674, -75.15059, -86.38568, -78.2986, 
    -89.73518, -78.6766, -92.43329, -78.98061, -90.99026, -79.30116, 
    -95.02118, -79.54681, -102.4268, -79.85341, -105.9435, -80.10781, -60, 
    -80.20015, -104.8801, -80.54588, -60, -80.72876, -101.5117, -80.92246, 
    -60, -81.00877, -60, -81.06235, -60, -81.1608, -106.4742, -81.29718, 
    -103.9641, -81.37227, -60, -81.3616, -60, -81.40285, _, _, _,
  37.88027, 37.86631, 37.87635, 37.86631, 37.88027, 37.88027, 37.87635, 
    37.86631, 37.88027, 37.88027, 37.87635, 37.88027, 37.88027, 37.86631, 
    34.69432, -26.64984, -63.67447, -51.64482, -53.95557, -60.68866, 
    -78.10041, -71.45501, -68.92828, -72.54437, -84.98619, -85.91365, 
    -76.88781, -79.19701, -89.73996, -86.84682, -81.1367, -83.18546, 
    -93.28663, -87.64732, -84.65588, -87.69238, -96.20338, -88.38165, 
    -85.27009, -88.29456, -60, -88.95349, -85.8811, -88.92185, -60, 
    -89.35487, -86.34439, -89.32329, -60, -89.71451, -86.67965, -89.65247, 
    -60, -90.07447, -86.97884, -89.95375, -60, -90.27973, -87.08813, 
    -90.19493, -112.6061, -90.3334, -87.25071, -90.36269, -60, -90.37988, 
    -87.33115, _, _,
  43.90087, 43.88691, 43.90087, 43.88691, 43.90087, 43.90087, 43.89695, 
    43.88691, 43.90087, 43.90087, 43.89695, 43.88691, 43.90087, 43.90087, 
    40.89057, -20.62926, -57.6539, -45.62382, -47.93489, -54.66795, 
    -72.07979, -65.43933, -62.90507, -66.52496, -78.96551, -79.8542, 
    -70.86678, -73.18546, -83.71949, -80.83016, -75.15059, -77.17548, 
    -87.27147, -81.61904, -78.63686, -79.59309, -90.18365, -82.35211, 
    -79.24456, -81.93767, -60, -83.00774, -79.83515, -82.86685, -60, 
    -83.34954, -80.29716, -83.2851, -60, -83.72718, -80.66069, -83.63617, 
    -60, -84.04095, -80.95227, -83.95191, -60, -84.25685, -81.04021, 
    -84.13803, -106.4742, -84.33965, -81.25626, -84.33166, -60, -84.36873, 
    -81.31423, -84.09198, _,
  37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 
    37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 37.88027, 
    37.88027, -44.91081, -59.44931, -66.13577, -70.54655, -73.83926, 
    -76.50502, -78.71399, -80.63277, -82.32097, -83.80496, -85.19013, 
    -86.45882, -87.51433, -88.61549, -89.73996, -91.94852, -91.61378, 
    -92.44866, -94.68334, -95.70703, -94.53887, -97.43819, -98.78764, 
    -96.61922, -60, -60, -60, -101.7445, -102.6123, -60, -111.9621, 
    -109.8821, -60, -106.33, -108.9633, -110.4342, -112.2896, -60, -60, 
    -109.6865, -60, -60, -60, -60, -60, -60, -60, -115.7018, -60, -60, -60, 
    -60, -60, -60 ;

 SpectralWidth =
  2.025983, 1.992853, 2.006343, 1.992853, 2.025983, 1.992853, 2.02595, 
    1.992853, 2.025983, 1.992853, 2.006343, 1.992853, 2.025983, 6.218236, 
    16.18475, 29.11437, 63.31838, 57.98458, 78.84911, 96.24792, 94.92109, 
    31.19421, 167.6288, 165.1624, 126.3155, 181.2471, 189.3386, 186.6803, 
    54.00056, 6.230806, 6.023754, 165.6705, 122.9799, 6.213971, 6.288617, 
    6.333627, 2.708325, 6.752519, 6.454357, 6.495016, 1.752841, 6.20906, 
    6.224329, 6.268034, 2.606797, 6.209067, 7.379832, 6.437248, 1.752841, 
    6.218138, 7.285558, 6.410694, 1.752841, 6.217628, 6.397143, 6.24549, 
    1.752841, 6.235815, 7.694444, 6.380661, _, _, _, _, _, _, _, _, _,
  1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 
    1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 4.250353, 
    17.07026, 27.05707, 34.61575, 41.67736, 46.61252, 52.28283, 57.8309, 
    61.84081, 63.45279, 65.94059, 70.38137, 69.34791, 71.39738, 68.27331, 
    76.83926, 81.91822, 31.34323, 36.97963, 77.39622, 75.75794, 81.93385, 
    1.079564, 1.079564, 17.84664, 1.079564, 22.785, 22.14141, 5.470537, 
    18.34183, 1.079564, 2.939651, 1.079564, 1.079564, 1.079564, 1.079564, 
    1.079564, 1.079564, 1.079564, 1.079564, 1.25187, 1.767322, 1.079564, 
    1.079564, 1.079564, 1.079564, 1.079564, 1.079564, _, _, _, _, _, _, _, _,
  2.025983, 2.025983, 2.025983, 2.025983, 2.025983, 2.025983, 2.025983, 
    2.025983, 2.025983, 2.025983, 2.025983, 2.025983, 2.025983, 6.901467, 
    27.7164, 43.93177, 56.20435, 67.66971, 75.68388, 84.88662, 93.90255, 
    100.4803, 102.962, 107.0645, 114.3457, 112.6065, 115.9278, 110.8448, 
    124.7708, 132.4257, 50.88874, 60.04976, 125.6682, 122.9799, 133.1309, 
    1.752841, 1.752841, 28.9818, 1.752841, 51.94084, 35.94864, 8.887363, 
    29.77874, 1.752841, 4.774203, 1.752841, 1.752841, 1.752841, 1.752841, 
    1.752841, 1.752841, 1.752841, 1.752841, 2.034461, 2.869539, 1.752841, 
    1.752841, 1.752841, 1.752841, 1.752841, 1.752841, 3.373617, _, _, _, _, 
    _, _, _,
  1.247791, 1.227386, 1.247774, 1.247777, 1.247791, 1.247779, 1.235695, 
    1.247776, 1.247791, 1.247777, 1.235695, 1.247782, 1.247791, 1.037671, 
    3.24881, 6.207905, 31.46173, 26.39258, 34.97684, 13.10279, 50.70974, 
    67.87524, 86.35033, 3.713161, 64.24362, 105.2504, 3.714536, 3.701796, 
    77.04771, 115.1805, 3.720505, 3.841109, 36.97963, 3.727749, 3.872986, 
    3.929565, 1.079564, 3.906224, 50.80981, 3.916715, 1.079564, 3.887054, 
    3.973067, 3.831341, 1.628666, 3.990041, 3.87196, 3.92597, 1.079564, 
    3.962504, 3.936933, 3.838386, 1.079564, 3.820977, 3.867725, 3.80345, 
    1.316583, 3.838906, 3.94682, 4.317171, 1.079564, 3.90783, 3.834519, _, _, 
    _, _, _, _,
  2.025983, 1.992853, 2.025956, 2.025961, 2.025983, 2.025961, 2.02595, 
    1.992853, 2.025983, 1.992853, 2.02595, 2.025966, 2.025983, 1.684821, 
    5.274932, 10.07949, 51.08475, 42.80785, 56.74717, 21.28427, 82.30781, 
    110.6204, 140.3486, 6.025659, 104.3075, 171.0231, 6.045039, 6.000047, 
    125.0914, 187.2558, 6.043629, 6.231971, 60.04976, 165.6705, 6.289675, 
    6.2306, 1.752841, 6.332061, 6.42939, 6.217153, 1.752841, 6.317334, 
    6.432657, 6.216043, 2.644717, 6.475397, 6.42447, 6.383591, 1.752841, 
    6.275231, 6.408667, 6.223674, 1.752841, 6.233538, 6.288871, 6.253023, 
    2.131801, 6.388801, 6.429002, 6.248552, 1.752841, 7.088287, 6.241844, 
    6.269206, _, _, _, _, _,
  1.247791, 1.247774, 1.247791, 1.247775, 1.247791, 1.247774, 1.247791, 
    1.235695, 1.247791, 1.235695, 1.247791, 1.235695, 1.247791, 1.247101, 
    6.049928, 5.051492, 27.05707, 20.55033, 40.8378, 39.21779, 52.70932, 
    63.92324, 58.49231, 19.14864, 69.06918, 3.730744, 71.58612, 3.717483, 
    29.65938, 115.2076, 73.36575, 3.720505, 31.34323, 3.711869, 22.48142, 
    3.877581, 86.24947, 3.86293, 24.50707, 3.853584, 1.531952, 3.956169, 
    2.651083, 3.962895, 1.079564, 3.967269, 1.878798, 3.953378, 1.079564, 
    3.93993, 1.177225, 3.840122, 1.079564, 3.844008, 1.079564, 4.359474, 
    1.079564, 3.863629, 1.239267, 3.94036, 1.096146, 3.930106, 1.079564, 
    3.836321, 1.079564, _, _, _, _,
  2.025983, 2.02595, 2.025983, 2.006343, 2.025983, 2.006343, 2.025983, 
    2.006343, 2.025983, 2.025958, 2.025983, 2.006343, 2.025983, 2.006343, 
    9.823023, 12.52936, 43.93177, 33.34898, 66.31935, 63.68274, 85.58031, 
    103.7043, 94.92109, 145.7891, 112.1536, 178.6143, 116.2304, 192.5571, 
    48.15004, 187.0675, 119.1158, 6.043629, 50.88874, 6.023754, 36.50131, 
    6.298687, 140.0641, 6.278718, 39.78637, 6.246871, 2.491961, 6.438747, 
    4.304021, 6.431386, 1.752841, 48.08473, 3.052284, 6.247384, 1.752841, 
    6.399056, 1.899956, 6.243686, 1.752841, 6.245381, 1.752841, 7.285558, 
    1.752841, 7.158381, 1.975737, 6.243136, 1.779246, 6.391057, 1.752841, 
    6.224598, 1.752841, 6.403839, _, _, _,
  1.247791, 1.227386, 1.235695, 1.227386, 1.247791, 1.247776, 1.235695, 
    1.227386, 1.247791, 1.247784, 1.235695, 1.247779, 1.247791, 1.227386, 
    1.079564, 3.543665, 22.42192, 8.412159, 23.75206, 33.51837, 49.64824, 
    14.97985, 67.3034, 73.61272, 63.7873, 3.709883, 110.6875, 106.9954, 
    68.70052, 3.690426, 115.2076, 115.1805, 81.91822, 3.832758, 3.7115, 
    3.73924, 71.69566, 3.831555, 3.871216, 3.88933, 1.079564, 3.908161, 
    3.966007, 3.887409, 1.079564, 3.819587, 3.854039, 3.877801, 1.079564, 
    3.902018, 3.918899, 3.931573, 1.079564, 3.828231, 3.948549, 3.962606, 
    1.079564, 3.848247, 3.920337, 3.911279, 1.239267, 3.936325, 3.94682, 
    3.851668, 1.079564, 3.931288, 4.832363, _, _,
  2.025983, 1.992853, 2.025956, 1.992853, 2.025983, 2.025967, 2.006343, 
    1.992853, 2.025983, 2.025965, 2.006343, 1.992853, 2.025983, 2.025878, 
    0.7152159, 5.75368, 36.40549, 13.65754, 38.55056, 54.28288, 80.6097, 
    24.30852, 109.4798, 119.596, 103.5706, 6.025446, 180.0124, 173.9689, 
    111.5496, 6.002167, 187.0675, 187.2558, 132.4257, 6.230806, 6.025172, 
    168.64, 116.4174, 6.21583, 6.291247, 23.88896, 1.752841, 6.368627, 
    6.448733, 6.31375, 1.752841, 6.206863, 6.413168, 6.274366, 1.752841, 
    6.224619, 6.392383, 6.46539, 1.752841, 6.209785, 6.402837, 6.425052, 
    1.752841, 6.232766, 6.356307, 6.466734, 1.975737, 6.401738, 6.429002, 
    6.257268, 1.752841, 6.372935, 7.694444, 6.338221, _,
  1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 
    1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 1.247791, 
    1.247791, 6.049928, 17.07026, 25.94239, 33.53618, 40.70324, 46.37259, 
    52.18637, 54.72458, 57.57774, 61.84081, 65.00509, 70.51196, 74.12808, 
    73.58384, 68.70052, 29.65938, 77.04771, 76.83926, 33.25862, 30.36143, 
    82.27775, 29.85907, 21.37081, 81.44975, 1.079564, 1.079564, 1.079564, 
    26.15518, 24.74459, 1.079564, 2.651083, 3.467576, 1.079564, 18.34183, 
    1.61655, 1.481648, 1.106439, 1.079564, 1.079564, 1.763889, 1.079564, 
    1.079564, 1.079564, 1.079564, 1.079564, 1.079564, 1.079564, 1.316583, 
    1.079564, 1.079564, 1.079564, 1.079564, 1.079564, 1.079564 ;

 NoiseLevel =
  -59.79054, -79.91229, -76.92703, -80.01283, -59.7893, -82.08401, -55.4295, 
    -83.50375, -59.79067, -91.09029, -87.4192, -90.05754, -62.81679, 
    -112.1676, -113.6862, -111.3251, -114.5785, -132.2387, -118.6768, 
    -115.3022, -117.2221, -119.0634, -123.019, -117.6744, -120.6432, 
    -132.9738, -125.8151, -120.9693, -117.7676, -125.4812, -113.1834, 
    -123.6707, -124.5995, -127.8893, -116.6471, -115.2313, -121.0981, 
    -134.7691, -120.235, -118.3479, -122.5352, -130.8357, -123.2721, 
    -120.4899, -124.8681, -130.9792, -137.1929, -123.0586, -126.426, 
    -130.1336, -138.0387, -125.2646, -128.0518, -129.6944, -128.9985, 
    -127.3342, -129.4005, -129.7838, -136.8324, -128.422, _, _, _, _, _, _, 
    _, _, _,
  -65.81114, -65.8102, -65.80978, -65.80941, -65.80951, -65.80969, -65.80991, 
    -65.81043, -65.81107, -65.81281, -65.81801, -65.84511, -66.38687, 
    -119.0371, -119.3562, -119.8634, -120.6682, -121.4972, -122.7696, 
    -122.2179, -123.2074, -124.7162, -126.3178, -125.2408, -126.5264, 
    -126.0039, -127.8265, -129.7301, -128.685, -129.384, -124.3949, 
    -125.4782, -130.3438, -130.6176, -134.9072, -127.032, -127.6891, 
    -128.0669, -127.9308, -128.8599, -130.4711, -129.6124, -130.386, 
    -129.9485, -130.5745, -130.0535, -131.4676, -131.744, -131.784, 
    -133.4083, -133.1307, -133.1049, -133.6704, -136.2254, -135.6491, 
    -135.6163, -135.6015, -134.8164, -135.3792, -135.9918, -135.8203, _, _, 
    _, _, _, _, _, _,
  -59.79054, -59.7896, -59.78918, -59.78881, -59.78891, -59.78909, -59.78931, 
    -59.78983, -59.79048, -59.79221, -59.79741, -59.82451, -60.36627, 
    -113.0763, -113.3397, -113.8436, -114.6477, -115.4763, -116.7469, 
    -116.1964, -117.1883, -118.7537, -120.2181, -119.2192, -120.5682, 
    -119.9864, -121.8038, -123.7024, -122.6632, -123.2909, -118.3695, 
    -119.4685, -124.3217, -124.5995, -129.0115, -120.9759, -121.6881, 
    -122.0345, -121.8643, -123.5479, -124.4604, -123.5841, -124.3697, 
    -123.9091, -124.5625, -124.0589, -125.4585, -125.6985, -125.7551, 
    -127.369, -127.0899, -127.0747, -127.5839, -130.2845, -129.6592, 
    -129.4194, -129.5396, -128.8227, -129.5993, -129.9493, -129.7411, 
    -128.848, _, _, _, _, _, _, _,
  -65.81114, -86.03049, -62.7135, -62.30402, -65.81023, -63.09006, -85.02598, 
    -61.63486, -65.81091, -62.33884, -92.4036, -69.01903, -65.9568, 
    -97.66461, -99.84877, -110.5166, -119.7559, -118.8036, -123.4239, 
    -118.9553, -122.1178, -121.8, -128.5532, -125.4663, -125.2253, -124.8677, 
    -117.3336, -126.7493, -127.9797, -128.3039, -117.8373, -131.2981, 
    -125.4782, -117.9958, -121.7662, -134.1552, -127.5577, -121.2593, 
    -142.4867, -136.4678, -127.941, -123.5641, -127.4967, -137.0059, 
    -128.9845, -126.5862, -130.2362, -136.562, -131.4416, -128.4534, 
    -132.6819, -136.8459, -134.2119, -130.9656, -134.2548, -136.223, 
    -135.4556, -132.6107, -135.4071, -144.3057, -134.4834, -133.9335, 
    -136.4387, _, _, _, _, _, _,
  -59.79054, -80.01857, -56.69289, -56.28336, -59.78962, -56.28508, 
    -55.42805, -86.10801, -59.79031, -86.21164, -55.71922, -60.2063, 
    -59.9362, -91.64146, -93.98022, -104.8446, -113.7386, -112.5682, 
    -116.7918, -113.1477, -116.0527, -115.759, -120.7344, -119.198, 
    -119.2046, -118.6488, -111.786, -120.4976, -121.954, -120.9328, 
    -111.3891, -124.9869, -119.4685, -123.6707, -115.2611, -128.219, 
    -121.5121, -114.9586, -118.7389, -129.2839, -121.9022, -117.4167, 
    -121.351, -130.1114, -122.9879, -120.4024, -123.7212, -130.3682, 
    -125.5292, -122.5519, -126.1824, -130.0702, -128.1834, -124.8543, 
    -128.1667, -129.7414, -129.3926, -126.788, -129.3746, -128.8652, 
    -128.4583, -133.2075, -130.2665, -128.8752, _, _, _, _, _,
  -65.81114, -62.70926, -65.81033, -63.2748, -65.80967, -62.72465, -65.81006, 
    -86.7508, -65.81062, -90.408, -65.81428, -93.4425, -65.86794, -65.98538, 
    -118.7152, -102.2059, -119.8634, -122.4245, -120.7445, -123.3017, 
    -123.1409, -125.8619, -123.2831, -114.9187, -125.8046, -117.4, -126.0569, 
    -117.4136, -121.8576, -134.6805, -129.7091, -117.8373, -124.3949, 
    -119.5193, -126.0421, -121.2646, -132.9309, -122.7127, -127.3546, 
    -124.1335, -126.4211, -126.1699, -129.2334, -127.1079, -128.5396, 
    -128.6941, -130.0023, -130.0132, -130.0535, -131.4017, -131.5255, 
    -132.0661, -132.2534, -133.1328, -133.0218, -144.9201, -133.5051, 
    -135.1537, -135.979, -135.8925, -145.3273, -135.8674, -134.4834, 
    -135.7369, -135.8203, _, _, _, _,
  -59.79054, -55.41281, -59.78974, -76.94506, -59.78907, -76.118, -59.78946, 
    -80.72209, -59.79002, -57.33859, -59.79368, -87.4192, -59.84734, 
    -90.3837, -112.6928, -113.4228, -113.8436, -115.2521, -114.728, 
    -116.8736, -117.1191, -119.1092, -117.2221, -121.4179, -119.7859, 
    -123.2639, -120.037, -126.7813, -115.8475, -127.811, -123.6846, 
    -111.3891, -118.3695, -113.1834, -120.0439, -115.1875, -126.9254, 
    -116.7058, -121.3762, -118.0546, -120.4067, -119.6007, -123.2032, 
    -120.885, -122.5352, -136.3775, -123.958, -123.7004, -124.0589, 
    -125.1968, -125.4802, -126.1189, -126.2336, -127.3117, -126.8993, 
    -138.0387, -127.5047, -137.3775, -129.8988, -129.3688, -139.1183, 
    -129.8325, -128.4583, -129.8166, -129.7411, -130.9241, _, _, _,
  -65.81114, -85.92162, -82.97549, -85.99834, -65.80988, -61.62906, 
    -84.09079, -87.73347, -65.81059, -67.02184, -91.50621, -63.38432, 
    -65.83863, -101.8705, -97.20427, -100.7556, -119.2318, -113.4223, 
    -122.0565, -118.8854, -122.57, -122.8737, -126.5037, -121.3513, 
    -124.4444, -126.4326, -130.9032, -125.1987, -127.1502, -126.5851, 
    -134.6805, -128.3039, -129.384, -131.3365, -119.5203, -118.055, 
    -133.4424, -134.1929, -122.3825, -120.9846, -127.3655, -135.6561, 
    -126.0439, -123.1406, -128.9755, -137.127, -128.2839, -126.1013, 
    -129.7284, -136.8326, -131.037, -127.6403, -131.1489, -136.2054, 
    -133.2083, -130.0754, -133.34, -137.27, -134.7322, -131.5871, -135.979, 
    -136.5883, -135.4071, -132.9914, -135.3792, -136.2929, -144.7204, _, _,
  -59.79054, -79.91199, -56.69223, -79.9953, -59.78927, -58.43605, -78.08126, 
    -81.71584, -59.78999, -57.73671, -85.47611, -88.1275, -59.81803, 
    -60.37433, -61.26431, -94.65394, -113.2111, -106.7014, -115.451, 
    -112.8373, -116.5473, -115.9123, -120.4573, -115.3284, -118.4225, 
    -121.0073, -123.1518, -118.8475, -121.1285, -120.4438, -127.811, 
    -120.9328, -123.2909, -125.4812, -113.1161, -124.1851, -127.4142, 
    -127.6938, -116.1447, -127.3836, -121.3653, -129.3498, -120.0542, 
    -116.8934, -122.9453, -130.6082, -122.1427, -119.6471, -123.6887, 
    -130.7983, -124.5722, -121.8247, -125.1247, -129.9526, -126.5325, 
    -124.037, -127.3087, -130.6971, -128.2381, -125.6135, -129.8988, 
    -130.3264, -129.3746, -126.7704, -129.5993, -129.8096, -136.8324, 
    -128.4741, _,
  -65.81114, -65.81036, -65.80998, -65.80991, -65.80977, -65.80989, 
    -65.80994, -65.81033, -65.81043, -65.81117, -65.81237, -65.81564, 
    -65.82587, -65.88662, -68.82005, -118.7152, -119.3562, -119.6891, 
    -120.8411, -121.178, -121.77, -122.7454, -123.2005, -122.9226, -124.7162, 
    -125.299, -125.431, -127.1485, -126.276, -127.1502, -121.8576, -127.9797, 
    -128.685, -123.7882, -123.9647, -131.085, -125.1177, -125.1628, 
    -132.2372, -126.6568, -127.032, -128.5842, -128.2324, -129.0974, 
    -127.0479, -129.2334, -129.4756, -128.4273, -130.386, -129.9989, 
    -130.0724, -129.6789, -130.6368, -131.4119, -131.765, -131.5265, 
    -133.4083, -133.3124, -133.34, -133.0634, -133.5051, -134.9247, 
    -135.4556, -135.2894, -135.6015, -135.6085, -135.3313, -135.5611, 
    -135.5345 ;
}
