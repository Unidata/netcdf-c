netcdf firstFile {
types:
  compound compoundType_3 {
    double member3(10) ;
  }; // compoundType_3
dimensions:
	dim3 = UNLIMITED ; // (1000 currently)
variables:
	compoundType_3 var_3(dim3) ;
		var_3:_Storage = "chunked" ;
		var_3:_ChunkSizes = 1000 ;
		var_3:_DeflateLevel = 1 ;
		var_3:_Shuffle = "true" ;
		//var_3:_Fletcher32 = "true" ;
		//var_3:_NoFill = "true" ;

// global attributes:
		:_Format = "netCDF-4" ;
data:

 var_3 = {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}}, 
    {{1, 2, 5, 10, 17, 0, 0, 0, 0, 0}} ;
}
