netcdf test_struct_nested {
types:
  compound x.field1_t {
    int x ;
    int y ;
  }; // x.field1_t
  compound x.field2_t {
    s1_t field1 ;
    s1_t field2 ;
  }; // x.field2_t
  compound x_t {
    x.field1_t field1 ;
    x.field1_t field2 ;
  }; // x_t
variables:
	x_t x ;
}
