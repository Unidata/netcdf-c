netcdf gfs.t00z.atmf024 {
dimensions:
	grid_xt = 3072 ;
	grid_yt = 1536 ;
	pfull = 127 ;
	phalf = 128 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:cartesian_axis = "X" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:units = "degrees_E" ;
		grid_xt:_Storage = "contiguous" ;
		grid_xt:_Endianness = "little" ;
	double lon(grid_yt, grid_xt) ;
		lon:long_name = "T-cell longitude" ;
		lon:units = "degrees_E" ;
		lon:_Storage = "contiguous" ;
		lon:_Endianness = "little" ;
	double grid_yt(grid_yt) ;
		grid_yt:cartesian_axis = "Y" ;
		grid_yt:long_name = "T-cell latiitude" ;
		grid_yt:units = "degrees_N" ;
		grid_yt:_Storage = "contiguous" ;
		grid_yt:_Endianness = "little" ;
	double lat(grid_yt, grid_xt) ;
		lat:long_name = "T-cell latitude" ;
		lat:units = "degrees_N" ;
		lat:_Storage = "contiguous" ;
		lat:_Endianness = "little" ;
	float pfull(pfull) ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:cartesian_axis = "Z" ;
		pfull:positive = "down" ;
		pfull:edges = "phalf" ;
		pfull:_Storage = "contiguous" ;
		pfull:_Endianness = "little" ;
	float phalf(phalf) ;
		phalf:long_name = "ref half pressure level" ;
		phalf:units = "mb" ;
		phalf:cartesian_axis = "Z" ;
		phalf:positive = "down" ;
		phalf:_Storage = "contiguous" ;
		phalf:_Endianness = "little" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "hours since 2018-01-10 00:00:00" ;
		time:cartesian_axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "JULIAN" ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 1 ;
		time:_Endianness = "little" ;
	float cld_amt(time, pfull, grid_yt, grid_xt) ;
		cld_amt:long_name = "cloud amount" ;
		cld_amt:units = "1" ;
		cld_amt:missing_value = -1.e+10f ;
		cld_amt:_FillValue = -1.e+10f ;
		cld_amt:cell_methods = "time: point" ;
		cld_amt:output_file = "atm" ;
		cld_amt:max_abs_compression_error = 3.057718e-05f ;
		cld_amt:nbits = 14 ;
		cld_amt:_Storage = "chunked" ;
		cld_amt:_ChunkSizes = 1, 22, 308, 615 ;
		cld_amt:_DeflateLevel = 1 ;
		cld_amt:_Endianness = "little" ;
	float clwmr(time, pfull, grid_yt, grid_xt) ;
		clwmr:long_name = "cloud water mixing ratio" ;
		clwmr:units = "kg/kg" ;
		clwmr:missing_value = -1.e+10f ;
		clwmr:_FillValue = -1.e+10f ;
		clwmr:cell_methods = "time: point" ;
		clwmr:output_file = "atm" ;
		clwmr:max_abs_compression_error = 4.976755e-08f ;
		clwmr:nbits = 14 ;
		clwmr:_Storage = "chunked" ;
		clwmr:_ChunkSizes = 1, 22, 308, 615 ;
		clwmr:_DeflateLevel = 1 ;
		clwmr:_Endianness = "little" ;
	float delz(time, pfull, grid_yt, grid_xt) ;
		delz:long_name = "height thickness" ;
		delz:units = "m" ;
		delz:missing_value = -1.e+10f ;
		delz:_FillValue = -1.e+10f ;
		delz:cell_methods = "time: point" ;
		delz:output_file = "atm" ;
		delz:max_abs_compression_error = 0.1002197f ;
		delz:nbits = 14 ;
		delz:_Storage = "chunked" ;
		delz:_ChunkSizes = 1, 22, 308, 615 ;
		delz:_DeflateLevel = 1 ;
		delz:_Endianness = "little" ;
	float dpres(time, pfull, grid_yt, grid_xt) ;
		dpres:long_name = "pressure thickness" ;
		dpres:units = "pa" ;
		dpres:missing_value = -1.e+10f ;
		dpres:_FillValue = -1.e+10f ;
		dpres:cell_methods = "time: point" ;
		dpres:output_file = "atm" ;
		dpres:max_abs_compression_error = 0.05603027f ;
		dpres:nbits = 14 ;
		dpres:_Storage = "chunked" ;
		dpres:_ChunkSizes = 1, 22, 308, 615 ;
		dpres:_DeflateLevel = 1 ;
		dpres:_Endianness = "little" ;
	float dzdt(time, pfull, grid_yt, grid_xt) ;
		dzdt:long_name = "vertical wind" ;
		dzdt:units = "m/sec" ;
		dzdt:missing_value = -1.e+10f ;
		dzdt:_FillValue = -1.e+10f ;
		dzdt:cell_methods = "time: point" ;
		dzdt:output_file = "atm" ;
		dzdt:max_abs_compression_error = 0.0003833771f ;
		dzdt:nbits = 14 ;
		dzdt:_Storage = "chunked" ;
		dzdt:_ChunkSizes = 1, 22, 308, 615 ;
		dzdt:_DeflateLevel = 1 ;
		dzdt:_Endianness = "little" ;
	float grle(time, pfull, grid_yt, grid_xt) ;
		grle:long_name = "graupel mixing ratio" ;
		grle:units = "kg/kg" ;
		grle:missing_value = -1.e+10f ;
		grle:_FillValue = -1.e+10f ;
		grle:cell_methods = "time: point" ;
		grle:output_file = "atm" ;
		grle:max_abs_compression_error = 3.105961e-07f ;
		grle:nbits = 14 ;
		grle:_Storage = "chunked" ;
		grle:_ChunkSizes = 1, 22, 308, 615 ;
		grle:_DeflateLevel = 1 ;
		grle:_Endianness = "little" ;
	float hgtsfc(time, grid_yt, grid_xt) ;
		hgtsfc:long_name = "surface geopotential height" ;
		hgtsfc:units = "gpm" ;
		hgtsfc:missing_value = -1.e+10f ;
		hgtsfc:_FillValue = -1.e+10f ;
		hgtsfc:cell_methods = "time: point" ;
		hgtsfc:output_file = "atm" ;
		hgtsfc:_Storage = "chunked" ;
		hgtsfc:_ChunkSizes = 1, 768, 1536 ;
		hgtsfc:_DeflateLevel = 1 ;
		hgtsfc:_Shuffle = "true" ;
		hgtsfc:_Endianness = "little" ;
	float icmr(time, pfull, grid_yt, grid_xt) ;
		icmr:long_name = "cloud ice mixing ratio" ;
		icmr:units = "kg/kg" ;
		icmr:missing_value = -1.e+10f ;
		icmr:_FillValue = -1.e+10f ;
		icmr:cell_methods = "time: point" ;
		icmr:output_file = "atm" ;
		icmr:max_abs_compression_error = 4.316098e-08f ;
		icmr:nbits = 14 ;
		icmr:_Storage = "chunked" ;
		icmr:_ChunkSizes = 1, 22, 308, 615 ;
		icmr:_DeflateLevel = 1 ;
		icmr:_Endianness = "little" ;
	float o3mr(time, pfull, grid_yt, grid_xt) ;
		o3mr:long_name = "ozone mixing ratio" ;
		o3mr:units = "kg/kg" ;
		o3mr:missing_value = -1.e+10f ;
		o3mr:_FillValue = -1.e+10f ;
		o3mr:cell_methods = "time: point" ;
		o3mr:output_file = "atm" ;
		o3mr:max_abs_compression_error = 5.438778e-10f ;
		o3mr:nbits = 14 ;
		o3mr:_Storage = "chunked" ;
		o3mr:_ChunkSizes = 1, 22, 308, 615 ;
		o3mr:_DeflateLevel = 1 ;
		o3mr:_Endianness = "little" ;
	float pressfc(time, grid_yt, grid_xt) ;
		pressfc:long_name = "surface pressure" ;
		pressfc:units = "pa" ;
		pressfc:missing_value = -1.e+10f ;
		pressfc:_FillValue = -1.e+10f ;
		pressfc:cell_methods = "time: point" ;
		pressfc:output_file = "atm" ;
		pressfc:_Storage = "chunked" ;
		pressfc:_ChunkSizes = 1, 768, 1536 ;
		pressfc:_DeflateLevel = 1 ;
		pressfc:_Shuffle = "true" ;
		pressfc:_Endianness = "little" ;
	float rwmr(time, pfull, grid_yt, grid_xt) ;
		rwmr:long_name = "rain mixing ratio" ;
		rwmr:units = "kg/kg" ;
		rwmr:missing_value = -1.e+10f ;
		rwmr:_FillValue = -1.e+10f ;
		rwmr:cell_methods = "time: point" ;
		rwmr:output_file = "atm" ;
		rwmr:max_abs_compression_error = 1.406297e-07f ;
		rwmr:nbits = 14 ;
		rwmr:_Storage = "chunked" ;
		rwmr:_ChunkSizes = 1, 22, 308, 615 ;
		rwmr:_DeflateLevel = 1 ;
		rwmr:_Endianness = "little" ;
	float snmr(time, pfull, grid_yt, grid_xt) ;
		snmr:long_name = "snow mixing ratio" ;
		snmr:units = "kg/kg" ;
		snmr:missing_value = -1.e+10f ;
		snmr:_FillValue = -1.e+10f ;
		snmr:cell_methods = "time: point" ;
		snmr:output_file = "atm" ;
		snmr:max_abs_compression_error = 6.280607e-08f ;
		snmr:nbits = 14 ;
		snmr:_Storage = "chunked" ;
		snmr:_ChunkSizes = 1, 22, 308, 615 ;
		snmr:_DeflateLevel = 1 ;
		snmr:_Endianness = "little" ;
	float spfh(time, pfull, grid_yt, grid_xt) ;
		spfh:long_name = "specific humidity" ;
		spfh:units = "kg/kg" ;
		spfh:missing_value = -1.e+10f ;
		spfh:_FillValue = -1.e+10f ;
		spfh:cell_methods = "time: point" ;
		spfh:output_file = "atm" ;
		spfh:max_abs_compression_error = 7.404014e-07f ;
		spfh:nbits = 14 ;
		spfh:_Storage = "chunked" ;
		spfh:_ChunkSizes = 1, 22, 308, 615 ;
		spfh:_DeflateLevel = 1 ;
		spfh:_Endianness = "little" ;
	float tmp(time, pfull, grid_yt, grid_xt) ;
		tmp:long_name = "temperature" ;
		tmp:units = "K" ;
		tmp:missing_value = -1.e+10f ;
		tmp:_FillValue = -1.e+10f ;
		tmp:cell_methods = "time: point" ;
		tmp:output_file = "atm" ;
		tmp:max_abs_compression_error = 0.004516602f ;
		tmp:nbits = 14 ;
		tmp:_Storage = "chunked" ;
		tmp:_ChunkSizes = 1, 22, 308, 615 ;
		tmp:_DeflateLevel = 1 ;
		tmp:_Endianness = "little" ;
	float ugrd(time, pfull, grid_yt, grid_xt) ;
		ugrd:long_name = "zonal wind" ;
		ugrd:units = "m/sec" ;
		ugrd:missing_value = -1.e+10f ;
		ugrd:_FillValue = -1.e+10f ;
		ugrd:cell_methods = "time: point" ;
		ugrd:output_file = "atm" ;
		ugrd:max_abs_compression_error = 0.008621216f ;
		ugrd:nbits = 14 ;
		ugrd:_Storage = "chunked" ;
		ugrd:_ChunkSizes = 1, 22, 308, 615 ;
		ugrd:_DeflateLevel = 1 ;
		ugrd:_Endianness = "little" ;
	float vgrd(time, pfull, grid_yt, grid_xt) ;
		vgrd:long_name = "meridional wind" ;
		vgrd:units = "m/sec" ;
		vgrd:missing_value = -1.e+10f ;
		vgrd:_FillValue = -1.e+10f ;
		vgrd:cell_methods = "time: point" ;
		vgrd:output_file = "atm" ;
		vgrd:max_abs_compression_error = 0.00667572f ;
		vgrd:nbits = 14 ;
		vgrd:_Storage = "chunked" ;
		vgrd:_ChunkSizes = 1, 22, 308, 615 ;
		vgrd:_DeflateLevel = 1 ;
		vgrd:_Endianness = "little" ;

// global attributes:
		:hydrostatic = "non-hydrostatic" ;
		:ncnsto = 9 ;
		:ak = 0.999f, 1.605f, 2.532f, 3.924f, 5.976f, 8.947f, 13.177f, 19.096f, 27.243f, 38.276f, 52.984f, 72.293f, 97.269f, 129.11f, 169.135f, 218.767f, 279.506f, 352.894f, 440.481f, 543.782f, 664.236f, 803.164f, 961.734f, 1140.931f, 1341.538f, 1564.119f, 1809.028f, 2076.415f, 2366.252f, 2678.372f, 3012.51f, 3368.363f, 3745.646f, 4144.164f, 4563.881f, 5004.995f, 5468.017f, 5953.848f, 6463.864f, 7000.f, 7563.494f, 8150.661f, 8756.529f, 9376.141f, 10004.55f, 10636.85f, 11268.16f, 11893.64f, 12508.52f, 13108.09f, 13687.73f, 14242.89f, 14769.15f, 15262.2f, 15717.86f, 16132.09f, 16501.02f, 16820.94f, 17088.32f, 17299.85f, 17453.08f, 17548.35f, 17586.77f, 17569.7f, 17498.7f, 17375.56f, 17202.3f, 16981.14f, 16714.5f, 16405.02f, 16055.49f, 15668.86f, 15248.25f, 14796.87f, 14318.04f, 13815.15f, 13291.63f, 12750.92f, 12196.47f, 11631.66f, 11059.83f, 10484.21f, 9907.927f, 9333.967f, 8765.155f, 8204.142f, 7653.387f, 7115.147f, 6591.468f, 6084.176f, 5594.876f, 5124.949f, 4675.554f, 4247.633f, 3841.918f, 3458.933f, 3099.01f, 2762.297f, 2448.768f, 2158.238f, 1890.375f, 1644.712f, 1420.661f, 1217.528f, 1034.524f, 870.778f, 725.348f, 597.235f, 485.392f, 388.734f, 306.149f, 236.502f, 178.651f, 131.447f, 93.74f, 64.392f, 42.274f, 26.274f, 15.302f, 8.287f, 4.19f, 1.994f, 0.81f, 0.232f, 0.029f, 0.f, 0.f, 0.f ;
		:bk = 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 1.018e-05f, 8.141e-05f, 0.00027469f, 0.00065078f, 0.00127009f, 0.00219248f, 0.00347713f, 0.00518228f, 0.00736504f, 0.0100812f, 0.01338492f, 0.01732857f, 0.02196239f, 0.02733428f, 0.03348954f, 0.04047056f, 0.04831661f, 0.05706358f, 0.06674372f, 0.07738548f, 0.08900629f, 0.101594f, 0.1151262f, 0.1295762f, 0.1449129f, 0.1611008f, 0.1780999f, 0.195866f, 0.2143511f, 0.2335031f, 0.2532663f, 0.2735822f, 0.294389f, 0.3156229f, 0.337218f, 0.3591072f, 0.3812224f, 0.4034951f, 0.4258572f, 0.4482413f, 0.4705813f, 0.492813f, 0.5148743f, 0.5367062f, 0.5582525f, 0.5794605f, 0.6002815f, 0.6206707f, 0.6405875f, 0.6599957f, 0.6788633f, 0.6971631f, 0.714872f, 0.7319713f, 0.7484465f, 0.7642871f, 0.7794867f, 0.7940422f, 0.8079541f, 0.8212263f, 0.8338652f, 0.8458801f, 0.8572826f, 0.8680866f, 0.8783077f, 0.8879632f, 0.8970718f, 0.9056532f, 0.9137284f, 0.9213187f, 0.9284464f, 0.9351338f, 0.9414037f, 0.9472789f, 0.9527821f, 0.957936f, 0.962763f, 0.9672851f, 0.971524f, 0.9755009f, 0.9792364f, 0.9827508f, 0.9860625f, 0.9891851f, 0.9921299f, 0.9949077f, 0.9975282f, 1.f ;
		:source = "FV3GFS" ;
		:grid = "gaussian" ;
		:im = 3072 ;
		:jm = 1536 ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 0 ;
		:_Format = "netCDF-4 classic model" ;
}
