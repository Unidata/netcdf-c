netcdf testmap {
dimensions:
	dim100 = 100 ;

group: _nczarr {
  } // group _nczarr

group: meta1 {

  // group attributes:
  		:data = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4]}" ;
  } // group meta1

group: meta2 {

  // group attributes:
  		:data = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4],\n\"extra\": 137}" ;
  } // group meta2

group: data1 {
  variables:
  	ubyte data(dim100) ;
  data:

   data = 0, 0, 0, 0, 1, 0, 0, 0, 2, 0, 0, 0, 3, 0, 0, 0, 4, 0, 0, 0, 5, 0, 
      0, 0, 6, 0, 0, 0, 7, 0, 0, 0, 8, 0, 0, 0, 9, 0, 0, 0, 10, 0, 0, 0, 11, 
      0, 0, 0, 12, 0, 0, 0, 13, 0, 0, 0, 14, 0, 0, 0, 15, 0, 0, 0, 16, 0, 0, 
      0, 17, 0, 0, 0, 18, 0, 0, 0, 19, 0, 0, 0, 20, 0, 0, 0, 21, 0, 0, 0, 22, 
      0, 0, 0, 23, 0, 0, 0, 24, 0, 0, 0 ;
  } // group data1
}
