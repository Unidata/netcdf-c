netcdf tmp_xarray {
dimensions:
	x = 2 ;
	y = 5 ;
variables:
	int i(x, y) ;
 		i:_FillValue = -2147483647 ;
data:

 i =
  _, _, _, _, _,
  _, _, _, _, _ ;
}
