netcdf ref_purezarr {
dimensions:
    x = 2;
    y = 5;
variables:
	int i(x,y) ;
}
