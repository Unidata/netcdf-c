netcdf testmap {

group: _nczarr {
  dimensions:
  	data_dim = UNLIMITED ; // (0 currently)
  variables:
  	ubyte data(data_dim) ;
  data:
  } // group _nczarr

group: meta1 {

  group: _zarray {
    dimensions:
    	data_dim = UNLIMITED ; // (50 currently)
    variables:
    	ubyte data(data_dim) ;
    data:

     data = 123, 10, 34, 102, 111, 111, 34, 58, 32, 52, 50, 44, 10, 34, 98, 
        97, 114, 34, 58, 32, 34, 97, 112, 112, 108, 101, 115, 34, 44, 10, 34, 
        98, 97, 122, 34, 58, 32, 91, 49, 44, 32, 50, 44, 32, 51, 44, 32, 52, 
        93, 125 ;
    } // group _zarray
  } // group meta1
}
