netcdf tmp_purezarr {
dimensions:
	_Anonymous_Dim_2 = 2 ;
	_Anonymous_Dim_5 = 5 ;
variables:
	int i(_Anonymous_Dim_2, _Anonymous_Dim_5) ;
	    i:_FillValue = -2147483647 ;
data:

 i =
  _, _, _, _, _,
  _, _, _, _, _ ;
}
