netcdf ref_any {
dimensions:
	dim0 = 4 ;
	dim1 = 4 ;
	dim2 = 4 ;
variables:
	int ivar(dim0, dim1, dim2) ;
 		ivar:_FillValue = -2147483647 ;
		ivar:_Storage = @chunked@ ;
		ivar:_ChunkSizes = 4, 4, 4 ;
		ivar:_Filter = @IH5@ ;
		ivar:_Codecs = @ICX@ ;
	float fvar(dim0, dim1, dim2) ;
 		fvar:_FillValue = 9.96921e+36f ;
		fvar:_Storage = @chunked@ ;
		fvar:_ChunkSizes = 4, 4, 4 ;
		fvar:_Filter = @FH5@ ;
		fvar:_Codecs = @FCX@ ;

data:

 ivar =
  0, 1, 2, 3,
  4, 5, 6, 7,
  8, 9, 10, 11,
  12, 13, 14, 15,
  16, 17, 18, 19,
  20, 21, 22, 23,
  24, 25, 26, 27,
  28, 29, 30, 31,
  32, 33, 34, 35,
  36, 37, 38, 39,
  40, 41, 42, 43,
  44, 45, 46, 47,
  48, 49, 50, 51,
  52, 53, 54, 55,
  56, 57, 58, 59,
  60, 61, 62, 63 ;

 fvar =
  0.5, 1.5, 2.5, 3.5,
  4.5, 5.5, 6.5, 7.5,
  8.5, 9.5, 10.5, 11.5,
  12.5, 13.5, 14.5, 15.5,
  16.5, 17.5, 18.5, 19.5,
  20.5, 21.5, 22.5, 23.5,
  24.5, 25.5, 26.5, 27.5,
  28.5, 29.5, 30.5, 31.5,
  32.5, 33.5, 34.5, 35.5,
  36.5, 37.5, 38.5, 39.5,
  40.5, 41.5, 42.5, 43.5,
  44.5, 45.5, 46.5, 47.5,
  48.5, 49.5, 50.5, 51.5,
  52.5, 53.5, 54.5, 55.5,
  56.5, 57.5, 58.5, 59.5,
  60.5, 61.5, 62.5, 63.5 ;
}
