netcdf nczarr2zarr {
dimensions:
	_zdim_8 = 8 ;
variables:
	int v(_zdim_8, _zdim_8) ;
		v:_FillValue = -1 ;
data:

 v =
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 1, 2, 3,
  _, _, _, _, 4, 5, 6, 7,
  _, _, _, _, 8, 9, 10, 11,
  _, _, _, _, 12, 13, 14, 15 ;
}
