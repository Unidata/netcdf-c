netcdf \2004050412_eta_211 {
dimensions:
	record = UNLIMITED ; // (1 currently)
	x = 135 ;
	y = 95 ;
	datetime_len = 21 ;
	nmodels = 1 ;
	ngrids = 1 ;
	nav = 1 ;
	nav_len = 100 ;
variables:
	double reftime(record) ;
		reftime:long_name = "reference time" ;
		reftime:units = "hours since 1992-1-1" ;
	double valtime(record) ;
		valtime:long_name = "valid time" ;
		valtime:units = "hours since 1992-1-1" ;
	char datetime(record, datetime_len) ;
		datetime:long_name = "reference date and time" ;
	float valtime_offset(record) ;
		valtime_offset:long_name = "hours from reference time" ;
		valtime_offset:units = "hours" ;
	int model_id(nmodels) ;
		model_id:long_name = "generating process ID number" ;
	char nav_model(nav, nav_len) ;
		nav_model:long_name = "navigation model name" ;
	int grid_type_code(nav) ;
		grid_type_code:long_name = "GRIB-1 GDS data representation type" ;
	char grid_type(nav, nav_len) ;
		grid_type:long_name = "GRIB-1 grid type" ;
	char grid_name(nav, nav_len) ;
		grid_name:long_name = "grid name" ;
	int grid_center(nav) ;
		grid_center:long_name = "GRIB-1 originating center ID" ;
	int grid_number(nav, ngrids) ;
		grid_number:long_name = "GRIB-1 catalogued grid numbers" ;
		grid_number:_FillValue = -9999 ;
	char x_dim(nav, nav_len) ;
		x_dim:long_name = "x dimension name" ;
	char y_dim(nav, nav_len) ;
		y_dim:long_name = "y dimension name" ;
	int Nx(nav) ;
		Nx:long_name = "number of points along x-axis" ;
	int Ny(nav) ;
		Ny:long_name = "number of points along y-axis" ;
	float La1(nav) ;
		La1:long_name = "latitude of first grid point" ;
		La1:units = "degrees_north" ;
	float Lo1(nav) ;
		Lo1:long_name = "longitude of first grid point" ;
		Lo1:units = "degrees_east" ;
	float Lov(nav) ;
		Lov:long_name = "orientation of the grid" ;
		Lov:units = "degrees_east" ;
	float Dx(nav) ;
		Dx:long_name = "x-direction grid length" ;
		Dx:units = "km" ;
	float Dy(nav) ;
		Dy:long_name = "y-direction grid length" ;
		Dy:units = "km" ;
	byte ProjFlag(nav) ;
		ProjFlag:long_name = "projection center flag" ;
	byte ResCompFlag(nav) ;
		ResCompFlag:long_name = "resolution and component flags" ;
	float Z_sfc(record, y, x) ;
		Z_sfc:long_name = "Geopotential height, gpm" ;
		Z_sfc:units = "gp m" ;
		Z_sfc:_FillValue = -9999.f ;
		Z_sfc:navigation = "nav" ;

// global attributes:
		:record = "reftime, valtime" ;
		:history = "2003-09-25 16:09:26 - created by gribtocdl 1.4 - 12.12.2002" ;
		:title = "CMC_reg_HGT_SFC_0_ps60km_2003092500_P000.grib" ;
		:Conventions = "NUWG" ;
		:version = 0. ;
}
