netcdf ref_fillonly {
dimensions:
	x = UNLIMITED ; // (6 currently)
variables:
	int i(x) ;
		i:_Storage = "chunked" ;
		i:_ChunkSizes = 6 ;
	float f(x) ;
		f:_FillValue = -9999.f ;
		f:_Storage = "chunked" ;
		f:_ChunkSizes = 6 ;

// global attributes:
		:_Format = "netCDF-4" ;
data:

 i = 1, 2, 3, 4, 5, 6 ;
}
