netcdf x3 {
dimensions:
	time = 10 ;
	lat = 2 ;
	lon = 4 ;
variables:
	float three_dmn_rec_var(time, lat, lon) ;
		three_dmn_rec_var:long_name = "three dimensional record variable" ;
		three_dmn_rec_var:units = "watt meter-2" ;
		three_dmn_rec_var:_FillValue = -99.f ;
data:

 three_dmn_rec_var =
  1, 2, 3, 4,
  5, 6, 7, 8,
  9, 10, 11, 12,
  13, 14, 15, 16,
  17, 18, 19, 20,
  21, 22, 23, 24,
  25, 26, 27, 28,
  29, 30, 31, 32,
  33, 34, 35, 36,
  37, 38, 39, 40,
  41, 42, 43, 44,
  45, 46, 47, 48,
  49, 50, 51, 52,
  53, 54, 55, 56,
  57, 58, 59, 60,
  61, 62, 63, 64,
  65, 66, 67, 68,
  69, 70, 71, 72,
  73, 74, 75, 76,
  77, 78, 79, 80 ;

}
