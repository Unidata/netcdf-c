netcdf tmp_whole {
dimensions:
	d0 = 8 ;
	d1 = 8 ;
variables:
	int v(d0, d1) ;
		v:_FillValue = -1 ;
data:

 v =
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 1, 2, 3,
  _, _, _, _, 4, 5, 6, 7,
  _, _, _, _, 8, 9, 10, 11,
  _, _, _, _, 12, 13, 14, 15 ;
}
