netcdf scope_ancestor_only {
types:
  ubyte enum test_enum_type {OPTION1 = 0, OPTION2 = 1, OPTION3 = 2} ;
dimensions:
  d1 = 1 ;
  d2 = 1 ;
group: test_group {
  variables:
  	test_enum_type test_variable(d1,d2) ;
  		test_enum_type test_variable:_FillValue = OPTION1 ;

  group: test_subgroup1 {

      group: test_subsubgroup {
      } // group test_subsubgroup

   } // group test_subgroup1

    group: test_subgroup2 {
    } // group test_subgroup2

  } // group test_group
}
