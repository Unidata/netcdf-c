netcdf type_preorder {

group: preorder {
types:
  ubyte enum test_enum_type {OPTION1 = 0, OPTION2 = 1, OPTION3 = 2} ;
} // group preorder

group: test_group {
  variables:
  	/preorder/test_enum_type test_variable ;
  		/preorder/test_enum_type test_variable:_FillValue = OPTION1 ;
  } // group test_group
}
