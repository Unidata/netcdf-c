netcdf ref_fixedstring {
dimensions:
	phony_dim_0 = 4 ;
variables:
	string v1 ;
	string vn(phony_dim_0) ;

// global attributes:
		:att1 = "abcd" ;
		string :attn = "abcd", "efgh", "ijkl", "mnop" ;
data:

 v1 = "abcd" ;

 vn = "abcd", "efgh", "ijkl", "mnop" ;
}
