netcdf keyword2 {
dimensions:
string = 128;
variables:
int string(string);
}
