netcdf tst_times_nc4 {
dimensions:
	time = 1 ;
	bnds = 2 ;
	t3 = UNLIMITED ; // (3 currently)
variables:
	double t1_days(time) ;
		t1_days:units = "days since 1500-1-1" ;
	double t1_days_case(time) ;
		t1_days_case:units = "DaYs since 1500-1-1" ;
	double t1_st_days(time) ;
		t1_st_days:calendar = "standard" ;
		t1_st_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_gr_days(time) ;
		t1_gr_days:calendar = "gregorian" ;
		t1_gr_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_pg_days(time) ;
		t1_pg_days:calendar = "proleptic_gregorian" ;
		t1_pg_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_nl_days(time) ;
		t1_nl_days:calendar = "noleap" ;
		t1_nl_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_365_days(time) ;
		t1_365_days:calendar = "365_day" ;
		t1_365_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_al_days(time) ;
		t1_al_days:calendar = "all_leap" ;
		t1_al_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_366_days(time) ;
		t1_366_days:calendar = "366_day" ;
		t1_366_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_360_days(time) ;
		t1_360_days:calendar = "360_day" ;
		t1_360_days:units = "days since 1500-01-01 00:00:00" ;
	double t1_jl_days(time) ;
		t1_jl_days:calendar = "julian" ;
		t1_jl_days:units = "days since 1500-01-01 00:00:00" ;
	double t2_days(time) ;
		string t2_days:units = "days since 2000-6-15 12:00" ;
	double t2_st_days(time) ;
		string t2_st_days:calendar = "standard" ;
		string t2_st_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_gr_days(time) ;
		string t2_gr_days:calendar = "gregorian" ;
		string t2_gr_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_pg_days(time) ;
		string t2_pg_days:calendar = "proleptic_gregorian" ;
		string t2_pg_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_pgt_days(time) ;
		string t2_pgt_days:calendar = "proleptic_gregorian" ;
		string t2_pgt_days:units = "days since 2000-06-15T12:00:00" ;
	double t2_nl_days(time) ;
		string t2_nl_days:calendar = "noleap" ;
		string t2_nl_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_365_days(time) ;
		string t2_365_days:calendar = "365_day" ;
		string t2_365_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_al_days(time) ;
		string t2_al_days:calendar = "all_leap" ;
		string t2_al_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_366_days(time) ;
		string t2_366_days:calendar = "366_day" ;
		string t2_366_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_360_days(time) ;
		string t2_360_days:calendar = "360_day" ;
		string t2_360_days:units = "days since 2000-06-15 12:00:00" ;
	double t2_jl_days(time) ;
		string t2_jl_days:calendar = "julian" ;
		string t2_jl_days:units = "days since 2000-06-15 12:00:00" ;
	int t3(t3) ;
		t3:units = "days since 1804-1-1" ;
		t3:calendar = "gregorian" ;
		t3:bounds = "t3_bnds" ;
		t3:time1 = 1 ; // "1804-01-02"
		t3:time2 = 5, 6 ; // "1804-01-06", "1804-01-07"
		t3:time3 = 7.125f, 8.75f ; // "1804-01-08 03", "1804-01-09 18"
		t3:time4 = 58.5, 59.5, 60.5 ;
		  // "1804-02-28 12", "1804-02-29 12", "1804-03-01 12"
		t3:time5 = 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120 ;
		  // "1804-04-10", "1804-04-11", "1804-04-12", "1804-04-13",
		  // "1804-04-14", "1804-04-15", "1804-04-16", "1804-04-17",
		  // "1804-04-18", "1804-04-19", "1804-04-20", "1804-04-21",
		  // "1804-04-22", "1804-04-23", "1804-04-24", "1804-04-25",
		  // "1804-04-26", "1804-04-27", "1804-04-28", "1804-04-29",
		  // "1804-04-30"
	double t3_bnds(t3, bnds) ;
	int t4 ;
		t4:units = "days" ;
		t4:att1 = 1 ;
		t4:att2 = 5, 6 ;
		t4:att3 = 7.125f, 8.75f ;
data:

 t1_days = "2009-01-01" ;

 t1_days_case = "2009-01-01" ;

 t1_st_days = "2009-01-01" ;

 t1_gr_days = "2009-01-01" ;

 t1_pg_days = "2009-01-01" ;

 t1_nl_days = "2009-01-01" ;

 t1_365_days = "2009-01-01" ;

 t1_al_days = "2009-01-01" ;

 t1_366_days = "2009-01-01" ;

 t1_360_days = "2009-01-01" ;

 t1_jl_days = "2009-01-01" ;

 t2_days = "2009-01-01" ;

 t2_st_days = "2009-01-01" ;

 t2_gr_days = "2009-01-01" ;

 t2_pg_days = "2009-01-01" ;

 t2_pgt_days = "2009-01-01" ;

 t2_nl_days = "2009-01-01" ;

 t2_365_days = "2009-01-01" ;

 t2_al_days = "2009-01-01" ;

 t2_366_days = "2009-01-01" ;

 t2_360_days = "2009-01-01" ;

 t2_jl_days = "2009-01-01" ;

 t3 = "1804-01-11", "1804-01-12", "1804-01-13" ;

 t3_bnds =
  "1804-01-10 12", "1804-01-11 12",
  "1804-01-11 12", "1804-01-12 12",
  "1804-01-12 12", "1804-01-13 12" ;

 t4 = _ ;
}
