netcdf testmapnc4 {

group: _nczarr {
  } // group _nczarr
}
