[0] /.zgroup : (0) ||
