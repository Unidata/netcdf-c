netcdf tst_mud4 {
dimensions:
	F0 = 1 ;
	F1 = 2 ;
	F2 = 3 ;
	F3 = 5 ;
	U0 = UNLIMITED ; // (1 currently)
	U1 = UNLIMITED ; // (2 currently)
	U2 = UNLIMITED ; // (3 currently)
	U3 = UNLIMITED ; // (5 currently)
variables:
	int ff(F1, F2) ;
		ff:_FillValue = -2147483647 ;
	int uf(U1, F2) ;
		uf:_FillValue = -2147483647 ;
	int fu(F1, U2) ;
		fu:_FillValue = -2147483647 ;
	int uu(U1, U2) ;
		uu:_FillValue = -2147483647 ;
	int ufff(U0, F1, F2, F3) ;
		ufff:_FillValue = -2147483647 ;
	int uffu(U0, F1, F2, U3) ;
		uffu:_FillValue = -2147483647 ;
	int ufuf(U0, F1, U2, F3) ;
		ufuf:_FillValue = -2147483647 ;
	int ufuu(U0, F1, U2, U3) ;
		ufuu:_FillValue = -2147483647 ;
	int uuff(U0, U1, F2, F3) ;
		uuff:_FillValue = -2147483647 ;
	int uufu(U0, U1, F2, U3) ;
		uufu:_FillValue = -2147483647 ;
	int uuuf(U0, U1, U2, F3) ;
		uuuf:_FillValue = -2147483647 ;
	int uuuu(U0, U1, U2, U3) ;
		uuuu:_FillValue = -2147483647 ;
	int ffff(F0, F1, F2, F3) ;
		ffff:_FillValue = -2147483647 ;
data:

 ff =
  // ff(0, 0-2)
    1, 2, 3,
  // ff(1, 0-2)
    4, 5, 6 ;

 uf =
  // uf(0, 0-2)
    1, 2, 3,
  // uf(1, 0-2)
    4, 5, 6 ;

 fu =
  {// fu(0, 0-2)
    1, 2, 3},
  {// fu(1, 0-2)
    4, 5, 6} ;

 uu =
  {// uu(0, 0-2)
    1, 2, 3},
  {// uu(1, 0-2)
    4, 5, 6} ;

 ufff =
  // ufff(0,0,0, 0-4)
    1, 2, 3, 4, 5,
  // ufff(0,0,1, 0-4)
    6, 7, 8, 9, 10,
  // ufff(0,0,2, 0-4)
    11, 12, 13, 14, 15,
  // ufff(0,1,0, 0-4)
    16, 17, 18, 19, 20,
  // ufff(0,1,1, 0-4)
    21, 22, 23, 24, 25,
  // ufff(0,1,2, 0-4)
    26, 27, 28, 29, 30 ;

 uffu =
  {// uffu(0,0,0, 0-4)
    1, 2, 3, 4, 5},
  {// uffu(0,0,1, 0-4)
    6, 7, 8, 9, 10},
  {// uffu(0,0,2, 0-4)
    11, 12, 13, 14, 15},
  {// uffu(0,1,0, 0-4)
    16, 17, 18, 19, 20},
  {// uffu(0,1,1, 0-4)
    21, 22, 23, 24, 25},
  {// uffu(0,1,2, 0-4)
    26, 27, 28, 29, 30} ;

 ufuf =
  {// ufuf(0,0,0, 0-4)
    1, 2, 3, 4, 5,
  // ufuf(0,0,1, 0-4)
    6, 7, 8, 9, 10,
  // ufuf(0,0,2, 0-4)
    11, 12, 13, 14, 15},
  {// ufuf(0,1,0, 0-4)
    16, 17, 18, 19, 20,
  // ufuf(0,1,1, 0-4)
    21, 22, 23, 24, 25,
  // ufuf(0,1,2, 0-4)
    26, 27, 28, 29, 30} ;

 ufuu =
  {{// ufuu(0,0,0, 0-4)
    1, 2, 3, 4, 5},
  {// ufuu(0,0,1, 0-4)
    6, 7, 8, 9, 10},
  {// ufuu(0,0,2, 0-4)
    11, 12, 13, 14, 15}},
  {{// ufuu(0,1,0, 0-4)
    16, 17, 18, 19, 20},
  {// ufuu(0,1,1, 0-4)
    21, 22, 23, 24, 25},
  {// ufuu(0,1,2, 0-4)
    26, 27, 28, 29, 30}} ;

 uuff =
  {// uuff(0,0,0, 0-4)
    1, 2, 3, 4, 5,
  // uuff(0,0,1, 0-4)
    6, 7, 8, 9, 10,
  // uuff(0,0,2, 0-4)
    11, 12, 13, 14, 15,
  // uuff(0,1,0, 0-4)
    16, 17, 18, 19, 20,
  // uuff(0,1,1, 0-4)
    21, 22, 23, 24, 25,
  // uuff(0,1,2, 0-4)
    26, 27, 28, 29, 30} ;

 uufu =
  {{// uufu(0,0,0, 0-4)
    1, 2, 3, 4, 5},
  {// uufu(0,0,1, 0-4)
    6, 7, 8, 9, 10},
  {// uufu(0,0,2, 0-4)
    11, 12, 13, 14, 15},
  {// uufu(0,1,0, 0-4)
    16, 17, 18, 19, 20},
  {// uufu(0,1,1, 0-4)
    21, 22, 23, 24, 25},
  {// uufu(0,1,2, 0-4)
    26, 27, 28, 29, 30}} ;

 uuuf =
  {{// uuuf(0,0,0, 0-4)
    1, 2, 3, 4, 5,
  // uuuf(0,0,1, 0-4)
    6, 7, 8, 9, 10,
  // uuuf(0,0,2, 0-4)
    11, 12, 13, 14, 15},
  {// uuuf(0,1,0, 0-4)
    16, 17, 18, 19, 20,
  // uuuf(0,1,1, 0-4)
    21, 22, 23, 24, 25,
  // uuuf(0,1,2, 0-4)
    26, 27, 28, 29, 30}} ;

 uuuu =
  {{{// uuuu(0,0,0, 0-4)
    1, 2, 3, 4, 5},
  {// uuuu(0,0,1, 0-4)
    6, 7, 8, 9, 10},
  {// uuuu(0,0,2, 0-4)
    11, 12, 13, 14, 15}},
  {{// uuuu(0,1,0, 0-4)
    16, 17, 18, 19, 20},
  {// uuuu(0,1,1, 0-4)
    21, 22, 23, 24, 25},
  {// uuuu(0,1,2, 0-4)
    26, 27, 28, 29, 30}}} ;

 ffff =
  // ffff(0,0,0, 0-4)
    1, 2, 3, 4, 5,
  // ffff(0,0,1, 0-4)
    6, 7, 8, 9, 10,
  // ffff(0,0,2, 0-4)
    11, 12, 13, 14, 15,
  // ffff(0,1,0, 0-4)
    16, 17, 18, 19, 20,
  // ffff(0,1,1, 0-4)
    21, 22, 23, 24, 25,
  // ffff(0,1,2, 0-4)
    26, 27, 28, 29, 30 ;
}
