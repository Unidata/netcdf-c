netcdf c0 {
dimensions:
	Dr = UNLIMITED ;
	D1 = 1 ;
	D2 = 2 ;
	D3 = 3 ;
//	U  = UNLIMITED;
variables:
	char c1(D1);
	char cr(Dr) ;
	char cr2(Dr, D2) ;
	char cr21(Dr, D2, D1) ;
	char cr33(Dr, D3, D3) ;
data:
 c1 = "";
 cr = "a","b" ;
 cr2 =  "@",  "D",  "H",  "L" ;
 cr21 =  "@",  "D",  "H",  "L" ;
 cr33 =  "1", "two",  "3",  "4",  "5",  "six" ;
}
